--   _______    __    ______     ______     _____    ________
--  |   ____|  |  |  |   _  \   |   _  \   / __  \  |___  ___|
--  |  |____   |  |  |  |_|  |  |  |_| /  | |  | |     |  |
--  |   ____|  |  |  |       |  |   _  \  | |  | |     |  |
--  |  |____   |  |  |  |\  \   |  |_| |  | |__| |     |  |
--  |_______|  |__|  |__| \__\  |______/   \_____/     |__|
--
-- Module: TABLE_COSINUS
-- But: Infere une ROM avec SINUS
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity TABLE_SINUS is Port ( 
	H       : in  STD_LOGIC;
	ANGLE   : in  STD_LOGIC_VECTOR(15 downto 0);
	SINUS   : out STD_LOGIC_VECTOR(15 downto 0);
	COSINUS : out STD_LOGIC_VECTOR(15 downto 0)
);
end TABLE_SINUS;

architecture Behavioral of TABLE_SINUS is
TYPE tableSinus is array(0 to ((360+90)*8-1)) of STD_LOGIC_VECTOR(11 downto 0);
SIGNAL TABLE : tableSinus := (
X"000", X"004", X"009", X"00D", X"012", X"016", X"01B", X"01F", X"024", X"028", 
X"02D", X"031", X"036", X"03A", X"03F", X"043", X"047", X"04C", X"050", X"055", 
X"059", X"05E", X"062", X"067", X"06B", X"070", X"074", X"079", X"07D", X"081", 
X"086", X"08A", X"08F", X"093", X"098", X"09C", X"0A1", X"0A5", X"0AA", X"0AE", 
X"0B2", X"0B7", X"0BB", X"0C0", X"0C4", X"0C9", X"0CD", X"0D2", X"0D6", X"0DB", 
X"0DF", X"0E3", X"0E8", X"0EC", X"0F1", X"0F5", X"0FA", X"0FE", X"102", X"107", 
X"10B", X"110", X"114", X"119", X"11D", X"121", X"126", X"12A", X"12F", X"133", 
X"138", X"13C", X"140", X"145", X"149", X"14E", X"152", X"156", X"15B", X"15F", 
X"164", X"168", X"16C", X"171", X"175", X"17A", X"17E", X"182", X"187", X"18B", 
X"190", X"194", X"198", X"19D", X"1A1", X"1A5", X"1AA", X"1AE", X"1B3", X"1B7", 
X"1BB", X"1C0", X"1C4", X"1C8", X"1CD", X"1D1", X"1D5", X"1DA", X"1DE", X"1E2", 
X"1E7", X"1EB", X"1EF", X"1F4", X"1F8", X"1FC", X"201", X"205", X"209", X"20E", 
X"212", X"216", X"21B", X"21F", X"223", X"228", X"22C", X"230", X"235", X"239", 
X"23D", X"241", X"246", X"24A", X"24E", X"253", X"257", X"25B", X"25F", X"264", 
X"268", X"26C", X"270", X"275", X"279", X"27D", X"281", X"286", X"28A", X"28E", 
X"292", X"297", X"29B", X"29F", X"2A3", X"2A7", X"2AC", X"2B0", X"2B4", X"2B8", 
X"2BC", X"2C1", X"2C5", X"2C9", X"2CD", X"2D1", X"2D6", X"2DA", X"2DE", X"2E2", 
X"2E6", X"2EA", X"2EF", X"2F3", X"2F7", X"2FB", X"2FF", X"303", X"307", X"30C", 
X"310", X"314", X"318", X"31C", X"320", X"324", X"328", X"32D", X"331", X"335", 
X"339", X"33D", X"341", X"345", X"349", X"34D", X"351", X"355", X"359", X"35D", 
X"362", X"366", X"36A", X"36E", X"372", X"376", X"37A", X"37E", X"382", X"386", 
X"38A", X"38E", X"392", X"396", X"39A", X"39E", X"3A2", X"3A6", X"3AA", X"3AE", 
X"3B2", X"3B6", X"3BA", X"3BE", X"3C1", X"3C5", X"3C9", X"3CD", X"3D1", X"3D5", 
X"3D9", X"3DD", X"3E1", X"3E5", X"3E9", X"3ED", X"3F0", X"3F4", X"3F8", X"3FC", 
X"400", X"404", X"408", X"40C", X"40F", X"413", X"417", X"41B", X"41F", X"423", 
X"426", X"42A", X"42E", X"432", X"436", X"439", X"43D", X"441", X"445", X"449", 
X"44C", X"450", X"454", X"458", X"45B", X"45F", X"463", X"467", X"46A", X"46E", 
X"472", X"476", X"479", X"47D", X"481", X"484", X"488", X"48C", X"48F", X"493", 
X"497", X"49A", X"49E", X"4A2", X"4A5", X"4A9", X"4AD", X"4B0", X"4B4", X"4B7", 
X"4BB", X"4BF", X"4C2", X"4C6", X"4C9", X"4CD", X"4D1", X"4D4", X"4D8", X"4DB", 
X"4DF", X"4E2", X"4E6", X"4E9", X"4ED", X"4F0", X"4F4", X"4F7", X"4FB", X"4FE", 
X"502", X"505", X"509", X"50C", X"510", X"513", X"517", X"51A", X"51E", X"521", 
X"524", X"528", X"52B", X"52F", X"532", X"535", X"539", X"53C", X"540", X"543", 
X"546", X"54A", X"54D", X"550", X"554", X"557", X"55A", X"55E", X"561", X"564", 
X"568", X"56B", X"56E", X"571", X"575", X"578", X"57B", X"57F", X"582", X"585", 
X"588", X"58B", X"58F", X"592", X"595", X"598", X"59B", X"59F", X"5A2", X"5A5", 
X"5A8", X"5AB", X"5AE", X"5B2", X"5B5", X"5B8", X"5BB", X"5BE", X"5C1", X"5C4", 
X"5C7", X"5CA", X"5CE", X"5D1", X"5D4", X"5D7", X"5DA", X"5DD", X"5E0", X"5E3", 
X"5E6", X"5E9", X"5EC", X"5EF", X"5F2", X"5F5", X"5F8", X"5FB", X"5FE", X"601", 
X"604", X"607", X"60A", X"60D", X"60F", X"612", X"615", X"618", X"61B", X"61E", 
X"621", X"624", X"627", X"629", X"62C", X"62F", X"632", X"635", X"638", X"63A", 
X"63D", X"640", X"643", X"646", X"648", X"64B", X"64E", X"651", X"653", X"656", 
X"659", X"65C", X"65E", X"661", X"664", X"666", X"669", X"66C", X"66E", X"671", 
X"674", X"676", X"679", X"67B", X"67E", X"681", X"683", X"686", X"688", X"68B", 
X"68E", X"690", X"693", X"695", X"698", X"69A", X"69D", X"69F", X"6A2", X"6A4", 
X"6A7", X"6A9", X"6AC", X"6AE", X"6B1", X"6B3", X"6B6", X"6B8", X"6BA", X"6BD", 
X"6BF", X"6C2", X"6C4", X"6C6", X"6C9", X"6CB", X"6CE", X"6D0", X"6D2", X"6D5", 
X"6D7", X"6D9", X"6DB", X"6DE", X"6E0", X"6E2", X"6E5", X"6E7", X"6E9", X"6EB", 
X"6EE", X"6F0", X"6F2", X"6F4", X"6F6", X"6F9", X"6FB", X"6FD", X"6FF", X"701", 
X"704", X"706", X"708", X"70A", X"70C", X"70E", X"710", X"712", X"714", X"717", 
X"719", X"71B", X"71D", X"71F", X"721", X"723", X"725", X"727", X"729", X"72B", 
X"72D", X"72F", X"731", X"733", X"735", X"737", X"738", X"73A", X"73C", X"73E", 
X"740", X"742", X"744", X"746", X"748", X"749", X"74B", X"74D", X"74F", X"751", 
X"753", X"754", X"756", X"758", X"75A", X"75B", X"75D", X"75F", X"761", X"762", 
X"764", X"766", X"768", X"769", X"76B", X"76D", X"76E", X"770", X"771", X"773", 
X"775", X"776", X"778", X"77A", X"77B", X"77D", X"77E", X"780", X"781", X"783", 
X"784", X"786", X"788", X"789", X"78B", X"78C", X"78D", X"78F", X"790", X"792", 
X"793", X"795", X"796", X"798", X"799", X"79A", X"79C", X"79D", X"79F", X"7A0", 
X"7A1", X"7A3", X"7A4", X"7A5", X"7A7", X"7A8", X"7A9", X"7AA", X"7AC", X"7AD", 
X"7AE", X"7AF", X"7B1", X"7B2", X"7B3", X"7B4", X"7B6", X"7B7", X"7B8", X"7B9", 
X"7BA", X"7BB", X"7BD", X"7BE", X"7BF", X"7C0", X"7C1", X"7C2", X"7C3", X"7C4", 
X"7C5", X"7C6", X"7C7", X"7C8", X"7C9", X"7CB", X"7CC", X"7CD", X"7CE", X"7CE", 
X"7CF", X"7D0", X"7D1", X"7D2", X"7D3", X"7D4", X"7D5", X"7D6", X"7D7", X"7D8", 
X"7D9", X"7DA", X"7DA", X"7DB", X"7DC", X"7DD", X"7DE", X"7DF", X"7DF", X"7E0", 
X"7E1", X"7E2", X"7E2", X"7E3", X"7E4", X"7E5", X"7E5", X"7E6", X"7E7", X"7E7", 
X"7E8", X"7E9", X"7EA", X"7EA", X"7EB", X"7EB", X"7EC", X"7ED", X"7ED", X"7EE", 
X"7EE", X"7EF", X"7F0", X"7F0", X"7F1", X"7F1", X"7F2", X"7F2", X"7F3", X"7F3", 
X"7F4", X"7F4", X"7F5", X"7F5", X"7F6", X"7F6", X"7F7", X"7F7", X"7F7", X"7F8", 
X"7F8", X"7F9", X"7F9", X"7F9", X"7FA", X"7FA", X"7FA", X"7FB", X"7FB", X"7FB", 
X"7FC", X"7FC", X"7FC", X"7FC", X"7FD", X"7FD", X"7FD", X"7FD", X"7FE", X"7FE", 
X"7FE", X"7FE", X"7FE", X"7FF", X"7FF", X"7FF", X"7FF", X"7FF", X"7FF", X"7FF", 
X"800", X"800", X"800", X"800", X"800", X"800", X"800", X"800", X"800", X"800", 
X"800", X"800", X"800", X"800", X"800", X"800", X"800", X"800", X"800", X"800", 
X"800", X"7FF", X"7FF", X"7FF", X"7FF", X"7FF", X"7FF", X"7FF", X"7FE", X"7FE", 
X"7FE", X"7FE", X"7FE", X"7FD", X"7FD", X"7FD", X"7FD", X"7FC", X"7FC", X"7FC", 
X"7FC", X"7FB", X"7FB", X"7FB", X"7FA", X"7FA", X"7FA", X"7F9", X"7F9", X"7F9", 
X"7F8", X"7F8", X"7F7", X"7F7", X"7F7", X"7F6", X"7F6", X"7F5", X"7F5", X"7F4", 
X"7F4", X"7F3", X"7F3", X"7F2", X"7F2", X"7F1", X"7F1", X"7F0", X"7F0", X"7EF", 
X"7EE", X"7EE", X"7ED", X"7ED", X"7EC", X"7EB", X"7EB", X"7EA", X"7EA", X"7E9", 
X"7E8", X"7E7", X"7E7", X"7E6", X"7E5", X"7E5", X"7E4", X"7E3", X"7E2", X"7E2", 
X"7E1", X"7E0", X"7DF", X"7DF", X"7DE", X"7DD", X"7DC", X"7DB", X"7DA", X"7DA", 
X"7D9", X"7D8", X"7D7", X"7D6", X"7D5", X"7D4", X"7D3", X"7D2", X"7D1", X"7D0", 
X"7CF", X"7CE", X"7CE", X"7CD", X"7CC", X"7CB", X"7C9", X"7C8", X"7C7", X"7C6", 
X"7C5", X"7C4", X"7C3", X"7C2", X"7C1", X"7C0", X"7BF", X"7BE", X"7BD", X"7BB", 
X"7BA", X"7B9", X"7B8", X"7B7", X"7B6", X"7B4", X"7B3", X"7B2", X"7B1", X"7AF", 
X"7AE", X"7AD", X"7AC", X"7AA", X"7A9", X"7A8", X"7A7", X"7A5", X"7A4", X"7A3", 
X"7A1", X"7A0", X"79F", X"79D", X"79C", X"79A", X"799", X"798", X"796", X"795", 
X"793", X"792", X"790", X"78F", X"78D", X"78C", X"78B", X"789", X"788", X"786", 
X"784", X"783", X"781", X"780", X"77E", X"77D", X"77B", X"77A", X"778", X"776", 
X"775", X"773", X"771", X"770", X"76E", X"76D", X"76B", X"769", X"768", X"766", 
X"764", X"762", X"761", X"75F", X"75D", X"75B", X"75A", X"758", X"756", X"754", 
X"753", X"751", X"74F", X"74D", X"74B", X"749", X"748", X"746", X"744", X"742", 
X"740", X"73E", X"73C", X"73A", X"738", X"737", X"735", X"733", X"731", X"72F", 
X"72D", X"72B", X"729", X"727", X"725", X"723", X"721", X"71F", X"71D", X"71B", 
X"719", X"717", X"714", X"712", X"710", X"70E", X"70C", X"70A", X"708", X"706", 
X"704", X"701", X"6FF", X"6FD", X"6FB", X"6F9", X"6F6", X"6F4", X"6F2", X"6F0", 
X"6EE", X"6EB", X"6E9", X"6E7", X"6E5", X"6E2", X"6E0", X"6DE", X"6DB", X"6D9", 
X"6D7", X"6D5", X"6D2", X"6D0", X"6CE", X"6CB", X"6C9", X"6C6", X"6C4", X"6C2", 
X"6BF", X"6BD", X"6BA", X"6B8", X"6B6", X"6B3", X"6B1", X"6AE", X"6AC", X"6A9", 
X"6A7", X"6A4", X"6A2", X"69F", X"69D", X"69A", X"698", X"695", X"693", X"690", 
X"68E", X"68B", X"688", X"686", X"683", X"681", X"67E", X"67B", X"679", X"676", 
X"674", X"671", X"66E", X"66C", X"669", X"666", X"664", X"661", X"65E", X"65C", 
X"659", X"656", X"653", X"651", X"64E", X"64B", X"648", X"646", X"643", X"640", 
X"63D", X"63A", X"638", X"635", X"632", X"62F", X"62C", X"629", X"627", X"624", 
X"621", X"61E", X"61B", X"618", X"615", X"612", X"60F", X"60D", X"60A", X"607", 
X"604", X"601", X"5FE", X"5FB", X"5F8", X"5F5", X"5F2", X"5EF", X"5EC", X"5E9", 
X"5E6", X"5E3", X"5E0", X"5DD", X"5DA", X"5D7", X"5D4", X"5D1", X"5CE", X"5CA", 
X"5C7", X"5C4", X"5C1", X"5BE", X"5BB", X"5B8", X"5B5", X"5B2", X"5AE", X"5AB", 
X"5A8", X"5A5", X"5A2", X"59F", X"59B", X"598", X"595", X"592", X"58F", X"58B", 
X"588", X"585", X"582", X"57F", X"57B", X"578", X"575", X"571", X"56E", X"56B", 
X"568", X"564", X"561", X"55E", X"55A", X"557", X"554", X"550", X"54D", X"54A", 
X"546", X"543", X"540", X"53C", X"539", X"535", X"532", X"52F", X"52B", X"528", 
X"524", X"521", X"51E", X"51A", X"517", X"513", X"510", X"50C", X"509", X"505", 
X"502", X"4FE", X"4FB", X"4F7", X"4F4", X"4F0", X"4ED", X"4E9", X"4E6", X"4E2", 
X"4DF", X"4DB", X"4D8", X"4D4", X"4D1", X"4CD", X"4C9", X"4C6", X"4C2", X"4BF", 
X"4BB", X"4B7", X"4B4", X"4B0", X"4AD", X"4A9", X"4A5", X"4A2", X"49E", X"49A", 
X"497", X"493", X"48F", X"48C", X"488", X"484", X"481", X"47D", X"479", X"476", 
X"472", X"46E", X"46A", X"467", X"463", X"45F", X"45B", X"458", X"454", X"450", 
X"44C", X"449", X"445", X"441", X"43D", X"439", X"436", X"432", X"42E", X"42A", 
X"426", X"423", X"41F", X"41B", X"417", X"413", X"40F", X"40C", X"408", X"404", 
X"400", X"3FC", X"3F8", X"3F4", X"3F0", X"3ED", X"3E9", X"3E5", X"3E1", X"3DD", 
X"3D9", X"3D5", X"3D1", X"3CD", X"3C9", X"3C5", X"3C1", X"3BE", X"3BA", X"3B6", 
X"3B2", X"3AE", X"3AA", X"3A6", X"3A2", X"39E", X"39A", X"396", X"392", X"38E", 
X"38A", X"386", X"382", X"37E", X"37A", X"376", X"372", X"36E", X"36A", X"366", 
X"362", X"35D", X"359", X"355", X"351", X"34D", X"349", X"345", X"341", X"33D", 
X"339", X"335", X"331", X"32D", X"328", X"324", X"320", X"31C", X"318", X"314", 
X"310", X"30C", X"307", X"303", X"2FF", X"2FB", X"2F7", X"2F3", X"2EF", X"2EA", 
X"2E6", X"2E2", X"2DE", X"2DA", X"2D6", X"2D1", X"2CD", X"2C9", X"2C5", X"2C1", 
X"2BC", X"2B8", X"2B4", X"2B0", X"2AC", X"2A7", X"2A3", X"29F", X"29B", X"297", 
X"292", X"28E", X"28A", X"286", X"281", X"27D", X"279", X"275", X"270", X"26C", 
X"268", X"264", X"25F", X"25B", X"257", X"253", X"24E", X"24A", X"246", X"241", 
X"23D", X"239", X"235", X"230", X"22C", X"228", X"223", X"21F", X"21B", X"216", 
X"212", X"20E", X"209", X"205", X"201", X"1FC", X"1F8", X"1F4", X"1EF", X"1EB", 
X"1E7", X"1E2", X"1DE", X"1DA", X"1D5", X"1D1", X"1CD", X"1C8", X"1C4", X"1C0", 
X"1BB", X"1B7", X"1B3", X"1AE", X"1AA", X"1A5", X"1A1", X"19D", X"198", X"194", 
X"190", X"18B", X"187", X"182", X"17E", X"17A", X"175", X"171", X"16C", X"168", 
X"164", X"15F", X"15B", X"156", X"152", X"14E", X"149", X"145", X"140", X"13C", 
X"138", X"133", X"12F", X"12A", X"126", X"121", X"11D", X"119", X"114", X"110", 
X"10B", X"107", X"102", X"0FE", X"0FA", X"0F5", X"0F1", X"0EC", X"0E8", X"0E3", 
X"0DF", X"0DB", X"0D6", X"0D2", X"0CD", X"0C9", X"0C4", X"0C0", X"0BB", X"0B7", 
X"0B2", X"0AE", X"0AA", X"0A5", X"0A1", X"09C", X"098", X"093", X"08F", X"08A", 
X"086", X"081", X"07D", X"079", X"074", X"070", X"06B", X"067", X"062", X"05E", 
X"059", X"055", X"050", X"04C", X"047", X"043", X"03F", X"03A", X"036", X"031", 
X"02D", X"028", X"024", X"01F", X"01B", X"016", X"012", X"00D", X"009", X"004", 
X"000", X"804", X"809", X"80D", X"812", X"816", X"81B", X"81F", X"824", X"828", 
X"82D", X"831", X"836", X"83A", X"83F", X"843", X"847", X"84C", X"850", X"855", 
X"859", X"85E", X"862", X"867", X"86B", X"870", X"874", X"879", X"87D", X"881", 
X"886", X"88A", X"88F", X"893", X"898", X"89C", X"8A1", X"8A5", X"8AA", X"8AE", 
X"8B2", X"8B7", X"8BB", X"8C0", X"8C4", X"8C9", X"8CD", X"8D2", X"8D6", X"8DB", 
X"8DF", X"8E3", X"8E8", X"8EC", X"8F1", X"8F5", X"8FA", X"8FE", X"902", X"907", 
X"90B", X"910", X"914", X"919", X"91D", X"921", X"926", X"92A", X"92F", X"933", 
X"938", X"93C", X"940", X"945", X"949", X"94E", X"952", X"956", X"95B", X"95F", 
X"964", X"968", X"96C", X"971", X"975", X"97A", X"97E", X"982", X"987", X"98B", 
X"990", X"994", X"998", X"99D", X"9A1", X"9A5", X"9AA", X"9AE", X"9B3", X"9B7", 
X"9BB", X"9C0", X"9C4", X"9C8", X"9CD", X"9D1", X"9D5", X"9DA", X"9DE", X"9E2", 
X"9E7", X"9EB", X"9EF", X"9F4", X"9F8", X"9FC", X"A01", X"A05", X"A09", X"A0E", 
X"A12", X"A16", X"A1B", X"A1F", X"A23", X"A28", X"A2C", X"A30", X"A35", X"A39", 
X"A3D", X"A41", X"A46", X"A4A", X"A4E", X"A53", X"A57", X"A5B", X"A5F", X"A64", 
X"A68", X"A6C", X"A70", X"A75", X"A79", X"A7D", X"A81", X"A86", X"A8A", X"A8E", 
X"A92", X"A97", X"A9B", X"A9F", X"AA3", X"AA7", X"AAC", X"AB0", X"AB4", X"AB8", 
X"ABC", X"AC1", X"AC5", X"AC9", X"ACD", X"AD1", X"AD6", X"ADA", X"ADE", X"AE2", 
X"AE6", X"AEA", X"AEF", X"AF3", X"AF7", X"AFB", X"AFF", X"B03", X"B07", X"B0C", 
X"B10", X"B14", X"B18", X"B1C", X"B20", X"B24", X"B28", X"B2D", X"B31", X"B35", 
X"B39", X"B3D", X"B41", X"B45", X"B49", X"B4D", X"B51", X"B55", X"B59", X"B5D", 
X"B62", X"B66", X"B6A", X"B6E", X"B72", X"B76", X"B7A", X"B7E", X"B82", X"B86", 
X"B8A", X"B8E", X"B92", X"B96", X"B9A", X"B9E", X"BA2", X"BA6", X"BAA", X"BAE", 
X"BB2", X"BB6", X"BBA", X"BBE", X"BC1", X"BC5", X"BC9", X"BCD", X"BD1", X"BD5", 
X"BD9", X"BDD", X"BE1", X"BE5", X"BE9", X"BED", X"BF0", X"BF4", X"BF8", X"BFC", 
X"C00", X"C04", X"C08", X"C0C", X"C0F", X"C13", X"C17", X"C1B", X"C1F", X"C23", 
X"C26", X"C2A", X"C2E", X"C32", X"C36", X"C39", X"C3D", X"C41", X"C45", X"C49", 
X"C4C", X"C50", X"C54", X"C58", X"C5B", X"C5F", X"C63", X"C67", X"C6A", X"C6E", 
X"C72", X"C76", X"C79", X"C7D", X"C81", X"C84", X"C88", X"C8C", X"C8F", X"C93", 
X"C97", X"C9A", X"C9E", X"CA2", X"CA5", X"CA9", X"CAD", X"CB0", X"CB4", X"CB7", 
X"CBB", X"CBF", X"CC2", X"CC6", X"CC9", X"CCD", X"CD1", X"CD4", X"CD8", X"CDB", 
X"CDF", X"CE2", X"CE6", X"CE9", X"CED", X"CF0", X"CF4", X"CF7", X"CFB", X"CFE", 
X"D02", X"D05", X"D09", X"D0C", X"D10", X"D13", X"D17", X"D1A", X"D1E", X"D21", 
X"D24", X"D28", X"D2B", X"D2F", X"D32", X"D35", X"D39", X"D3C", X"D40", X"D43", 
X"D46", X"D4A", X"D4D", X"D50", X"D54", X"D57", X"D5A", X"D5E", X"D61", X"D64", 
X"D68", X"D6B", X"D6E", X"D71", X"D75", X"D78", X"D7B", X"D7F", X"D82", X"D85", 
X"D88", X"D8B", X"D8F", X"D92", X"D95", X"D98", X"D9B", X"D9F", X"DA2", X"DA5", 
X"DA8", X"DAB", X"DAE", X"DB2", X"DB5", X"DB8", X"DBB", X"DBE", X"DC1", X"DC4", 
X"DC7", X"DCA", X"DCE", X"DD1", X"DD4", X"DD7", X"DDA", X"DDD", X"DE0", X"DE3", 
X"DE6", X"DE9", X"DEC", X"DEF", X"DF2", X"DF5", X"DF8", X"DFB", X"DFE", X"E01", 
X"E04", X"E07", X"E0A", X"E0D", X"E0F", X"E12", X"E15", X"E18", X"E1B", X"E1E", 
X"E21", X"E24", X"E27", X"E29", X"E2C", X"E2F", X"E32", X"E35", X"E38", X"E3A", 
X"E3D", X"E40", X"E43", X"E46", X"E48", X"E4B", X"E4E", X"E51", X"E53", X"E56", 
X"E59", X"E5C", X"E5E", X"E61", X"E64", X"E66", X"E69", X"E6C", X"E6E", X"E71", 
X"E74", X"E76", X"E79", X"E7B", X"E7E", X"E81", X"E83", X"E86", X"E88", X"E8B", 
X"E8E", X"E90", X"E93", X"E95", X"E98", X"E9A", X"E9D", X"E9F", X"EA2", X"EA4", 
X"EA7", X"EA9", X"EAC", X"EAE", X"EB1", X"EB3", X"EB6", X"EB8", X"EBA", X"EBD", 
X"EBF", X"EC2", X"EC4", X"EC6", X"EC9", X"ECB", X"ECE", X"ED0", X"ED2", X"ED5", 
X"ED7", X"ED9", X"EDB", X"EDE", X"EE0", X"EE2", X"EE5", X"EE7", X"EE9", X"EEB", 
X"EEE", X"EF0", X"EF2", X"EF4", X"EF6", X"EF9", X"EFB", X"EFD", X"EFF", X"F01", 
X"F04", X"F06", X"F08", X"F0A", X"F0C", X"F0E", X"F10", X"F12", X"F14", X"F17", 
X"F19", X"F1B", X"F1D", X"F1F", X"F21", X"F23", X"F25", X"F27", X"F29", X"F2B", 
X"F2D", X"F2F", X"F31", X"F33", X"F35", X"F37", X"F38", X"F3A", X"F3C", X"F3E", 
X"F40", X"F42", X"F44", X"F46", X"F48", X"F49", X"F4B", X"F4D", X"F4F", X"F51", 
X"F53", X"F54", X"F56", X"F58", X"F5A", X"F5B", X"F5D", X"F5F", X"F61", X"F62", 
X"F64", X"F66", X"F68", X"F69", X"F6B", X"F6D", X"F6E", X"F70", X"F71", X"F73", 
X"F75", X"F76", X"F78", X"F7A", X"F7B", X"F7D", X"F7E", X"F80", X"F81", X"F83", 
X"F84", X"F86", X"F88", X"F89", X"F8B", X"F8C", X"F8D", X"F8F", X"F90", X"F92", 
X"F93", X"F95", X"F96", X"F98", X"F99", X"F9A", X"F9C", X"F9D", X"F9F", X"FA0", 
X"FA1", X"FA3", X"FA4", X"FA5", X"FA7", X"FA8", X"FA9", X"FAA", X"FAC", X"FAD", 
X"FAE", X"FAF", X"FB1", X"FB2", X"FB3", X"FB4", X"FB6", X"FB7", X"FB8", X"FB9", 
X"FBA", X"FBB", X"FBD", X"FBE", X"FBF", X"FC0", X"FC1", X"FC2", X"FC3", X"FC4", 
X"FC5", X"FC6", X"FC7", X"FC8", X"FC9", X"FCB", X"FCC", X"FCD", X"FCE", X"FCE", 
X"FCF", X"FD0", X"FD1", X"FD2", X"FD3", X"FD4", X"FD5", X"FD6", X"FD7", X"FD8", 
X"FD9", X"FDA", X"FDA", X"FDB", X"FDC", X"FDD", X"FDE", X"FDF", X"FDF", X"FE0", 
X"FE1", X"FE2", X"FE2", X"FE3", X"FE4", X"FE5", X"FE5", X"FE6", X"FE7", X"FE7", 
X"FE8", X"FE9", X"FEA", X"FEA", X"FEB", X"FEB", X"FEC", X"FED", X"FED", X"FEE", 
X"FEE", X"FEF", X"FF0", X"FF0", X"FF1", X"FF1", X"FF2", X"FF2", X"FF3", X"FF3", 
X"FF4", X"FF4", X"FF5", X"FF5", X"FF6", X"FF6", X"FF7", X"FF7", X"FF7", X"FF8", 
X"FF8", X"FF9", X"FF9", X"FF9", X"FFA", X"FFA", X"FFA", X"FFB", X"FFB", X"FFB", 
X"FFC", X"FFC", X"FFC", X"FFC", X"FFD", X"FFD", X"FFD", X"FFD", X"FFE", X"FFE", 
X"FFE", X"FFE", X"FFE", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", 
X"800", X"800", X"800", X"800", X"800", X"800", X"800", X"800", X"800", X"800", 
X"800", X"800", X"800", X"800", X"800", X"800", X"800", X"800", X"800", X"800", 
X"800", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFF", X"FFE", X"FFE", 
X"FFE", X"FFE", X"FFE", X"FFD", X"FFD", X"FFD", X"FFD", X"FFC", X"FFC", X"FFC", 
X"FFC", X"FFB", X"FFB", X"FFB", X"FFA", X"FFA", X"FFA", X"FF9", X"FF9", X"FF9", 
X"FF8", X"FF8", X"FF7", X"FF7", X"FF7", X"FF6", X"FF6", X"FF5", X"FF5", X"FF4", 
X"FF4", X"FF3", X"FF3", X"FF2", X"FF2", X"FF1", X"FF1", X"FF0", X"FF0", X"FEF", 
X"FEE", X"FEE", X"FED", X"FED", X"FEC", X"FEB", X"FEB", X"FEA", X"FEA", X"FE9", 
X"FE8", X"FE7", X"FE7", X"FE6", X"FE5", X"FE5", X"FE4", X"FE3", X"FE2", X"FE2", 
X"FE1", X"FE0", X"FDF", X"FDF", X"FDE", X"FDD", X"FDC", X"FDB", X"FDA", X"FDA", 
X"FD9", X"FD8", X"FD7", X"FD6", X"FD5", X"FD4", X"FD3", X"FD2", X"FD1", X"FD0", 
X"FCF", X"FCE", X"FCE", X"FCD", X"FCC", X"FCB", X"FC9", X"FC8", X"FC7", X"FC6", 
X"FC5", X"FC4", X"FC3", X"FC2", X"FC1", X"FC0", X"FBF", X"FBE", X"FBD", X"FBB", 
X"FBA", X"FB9", X"FB8", X"FB7", X"FB6", X"FB4", X"FB3", X"FB2", X"FB1", X"FAF", 
X"FAE", X"FAD", X"FAC", X"FAA", X"FA9", X"FA8", X"FA7", X"FA5", X"FA4", X"FA3", 
X"FA1", X"FA0", X"F9F", X"F9D", X"F9C", X"F9A", X"F99", X"F98", X"F96", X"F95", 
X"F93", X"F92", X"F90", X"F8F", X"F8D", X"F8C", X"F8B", X"F89", X"F88", X"F86", 
X"F84", X"F83", X"F81", X"F80", X"F7E", X"F7D", X"F7B", X"F7A", X"F78", X"F76", 
X"F75", X"F73", X"F71", X"F70", X"F6E", X"F6D", X"F6B", X"F69", X"F68", X"F66", 
X"F64", X"F62", X"F61", X"F5F", X"F5D", X"F5B", X"F5A", X"F58", X"F56", X"F54", 
X"F53", X"F51", X"F4F", X"F4D", X"F4B", X"F49", X"F48", X"F46", X"F44", X"F42", 
X"F40", X"F3E", X"F3C", X"F3A", X"F38", X"F37", X"F35", X"F33", X"F31", X"F2F", 
X"F2D", X"F2B", X"F29", X"F27", X"F25", X"F23", X"F21", X"F1F", X"F1D", X"F1B", 
X"F19", X"F17", X"F14", X"F12", X"F10", X"F0E", X"F0C", X"F0A", X"F08", X"F06", 
X"F04", X"F01", X"EFF", X"EFD", X"EFB", X"EF9", X"EF6", X"EF4", X"EF2", X"EF0", 
X"EEE", X"EEB", X"EE9", X"EE7", X"EE5", X"EE2", X"EE0", X"EDE", X"EDB", X"ED9", 
X"ED7", X"ED5", X"ED2", X"ED0", X"ECE", X"ECB", X"EC9", X"EC6", X"EC4", X"EC2", 
X"EBF", X"EBD", X"EBA", X"EB8", X"EB6", X"EB3", X"EB1", X"EAE", X"EAC", X"EA9", 
X"EA7", X"EA4", X"EA2", X"E9F", X"E9D", X"E9A", X"E98", X"E95", X"E93", X"E90", 
X"E8E", X"E8B", X"E88", X"E86", X"E83", X"E81", X"E7E", X"E7B", X"E79", X"E76", 
X"E74", X"E71", X"E6E", X"E6C", X"E69", X"E66", X"E64", X"E61", X"E5E", X"E5C", 
X"E59", X"E56", X"E53", X"E51", X"E4E", X"E4B", X"E48", X"E46", X"E43", X"E40", 
X"E3D", X"E3A", X"E38", X"E35", X"E32", X"E2F", X"E2C", X"E29", X"E27", X"E24", 
X"E21", X"E1E", X"E1B", X"E18", X"E15", X"E12", X"E0F", X"E0D", X"E0A", X"E07", 
X"E04", X"E01", X"DFE", X"DFB", X"DF8", X"DF5", X"DF2", X"DEF", X"DEC", X"DE9", 
X"DE6", X"DE3", X"DE0", X"DDD", X"DDA", X"DD7", X"DD4", X"DD1", X"DCE", X"DCA", 
X"DC7", X"DC4", X"DC1", X"DBE", X"DBB", X"DB8", X"DB5", X"DB2", X"DAE", X"DAB", 
X"DA8", X"DA5", X"DA2", X"D9F", X"D9B", X"D98", X"D95", X"D92", X"D8F", X"D8B", 
X"D88", X"D85", X"D82", X"D7F", X"D7B", X"D78", X"D75", X"D71", X"D6E", X"D6B", 
X"D68", X"D64", X"D61", X"D5E", X"D5A", X"D57", X"D54", X"D50", X"D4D", X"D4A", 
X"D46", X"D43", X"D40", X"D3C", X"D39", X"D35", X"D32", X"D2F", X"D2B", X"D28", 
X"D24", X"D21", X"D1E", X"D1A", X"D17", X"D13", X"D10", X"D0C", X"D09", X"D05", 
X"D02", X"CFE", X"CFB", X"CF7", X"CF4", X"CF0", X"CED", X"CE9", X"CE6", X"CE2", 
X"CDF", X"CDB", X"CD8", X"CD4", X"CD1", X"CCD", X"CC9", X"CC6", X"CC2", X"CBF", 
X"CBB", X"CB7", X"CB4", X"CB0", X"CAD", X"CA9", X"CA5", X"CA2", X"C9E", X"C9A", 
X"C97", X"C93", X"C8F", X"C8C", X"C88", X"C84", X"C81", X"C7D", X"C79", X"C76", 
X"C72", X"C6E", X"C6A", X"C67", X"C63", X"C5F", X"C5B", X"C58", X"C54", X"C50", 
X"C4C", X"C49", X"C45", X"C41", X"C3D", X"C39", X"C36", X"C32", X"C2E", X"C2A", 
X"C26", X"C23", X"C1F", X"C1B", X"C17", X"C13", X"C0F", X"C0C", X"C08", X"C04", 
X"C00", X"BFC", X"BF8", X"BF4", X"BF0", X"BED", X"BE9", X"BE5", X"BE1", X"BDD", 
X"BD9", X"BD5", X"BD1", X"BCD", X"BC9", X"BC5", X"BC1", X"BBE", X"BBA", X"BB6", 
X"BB2", X"BAE", X"BAA", X"BA6", X"BA2", X"B9E", X"B9A", X"B96", X"B92", X"B8E", 
X"B8A", X"B86", X"B82", X"B7E", X"B7A", X"B76", X"B72", X"B6E", X"B6A", X"B66", 
X"B62", X"B5D", X"B59", X"B55", X"B51", X"B4D", X"B49", X"B45", X"B41", X"B3D", 
X"B39", X"B35", X"B31", X"B2D", X"B28", X"B24", X"B20", X"B1C", X"B18", X"B14", 
X"B10", X"B0C", X"B07", X"B03", X"AFF", X"AFB", X"AF7", X"AF3", X"AEF", X"AEA", 
X"AE6", X"AE2", X"ADE", X"ADA", X"AD6", X"AD1", X"ACD", X"AC9", X"AC5", X"AC1", 
X"ABC", X"AB8", X"AB4", X"AB0", X"AAC", X"AA7", X"AA3", X"A9F", X"A9B", X"A97", 
X"A92", X"A8E", X"A8A", X"A86", X"A81", X"A7D", X"A79", X"A75", X"A70", X"A6C", 
X"A68", X"A64", X"A5F", X"A5B", X"A57", X"A53", X"A4E", X"A4A", X"A46", X"A41", 
X"A3D", X"A39", X"A35", X"A30", X"A2C", X"A28", X"A23", X"A1F", X"A1B", X"A16", 
X"A12", X"A0E", X"A09", X"A05", X"A01", X"9FC", X"9F8", X"9F4", X"9EF", X"9EB", 
X"9E7", X"9E2", X"9DE", X"9DA", X"9D5", X"9D1", X"9CD", X"9C8", X"9C4", X"9C0", 
X"9BB", X"9B7", X"9B3", X"9AE", X"9AA", X"9A5", X"9A1", X"99D", X"998", X"994", 
X"990", X"98B", X"987", X"982", X"97E", X"97A", X"975", X"971", X"96C", X"968", 
X"964", X"95F", X"95B", X"956", X"952", X"94E", X"949", X"945", X"940", X"93C", 
X"938", X"933", X"92F", X"92A", X"926", X"921", X"91D", X"919", X"914", X"910", 
X"90B", X"907", X"902", X"8FE", X"8FA", X"8F5", X"8F1", X"8EC", X"8E8", X"8E3", 
X"8DF", X"8DB", X"8D6", X"8D2", X"8CD", X"8C9", X"8C4", X"8C0", X"8BB", X"8B7", 
X"8B2", X"8AE", X"8AA", X"8A5", X"8A1", X"89C", X"898", X"893", X"88F", X"88A", 
X"886", X"881", X"87D", X"879", X"874", X"870", X"86B", X"867", X"862", X"85E", 
X"859", X"855", X"850", X"84C", X"847", X"843", X"83F", X"83A", X"836", X"831", 
X"82D", X"828", X"824", X"81F", X"81B", X"816", X"812", X"80D", X"809", X"804", 
X"000", X"004", X"009", X"00D", X"012", X"016", X"01B", X"01F", X"024", X"028", 
X"02D", X"031", X"036", X"03A", X"03F", X"043", X"047", X"04C", X"050", X"055", 
X"059", X"05E", X"062", X"067", X"06B", X"070", X"074", X"079", X"07D", X"081", 
X"086", X"08A", X"08F", X"093", X"098", X"09C", X"0A1", X"0A5", X"0AA", X"0AE", 
X"0B2", X"0B7", X"0BB", X"0C0", X"0C4", X"0C9", X"0CD", X"0D2", X"0D6", X"0DB", 
X"0DF", X"0E3", X"0E8", X"0EC", X"0F1", X"0F5", X"0FA", X"0FE", X"102", X"107", 
X"10B", X"110", X"114", X"119", X"11D", X"121", X"126", X"12A", X"12F", X"133", 
X"138", X"13C", X"140", X"145", X"149", X"14E", X"152", X"156", X"15B", X"15F", 
X"164", X"168", X"16C", X"171", X"175", X"17A", X"17E", X"182", X"187", X"18B", 
X"190", X"194", X"198", X"19D", X"1A1", X"1A5", X"1AA", X"1AE", X"1B3", X"1B7", 
X"1BB", X"1C0", X"1C4", X"1C8", X"1CD", X"1D1", X"1D5", X"1DA", X"1DE", X"1E2", 
X"1E7", X"1EB", X"1EF", X"1F4", X"1F8", X"1FC", X"201", X"205", X"209", X"20E", 
X"212", X"216", X"21B", X"21F", X"223", X"228", X"22C", X"230", X"235", X"239", 
X"23D", X"241", X"246", X"24A", X"24E", X"253", X"257", X"25B", X"25F", X"264", 
X"268", X"26C", X"270", X"275", X"279", X"27D", X"281", X"286", X"28A", X"28E", 
X"292", X"297", X"29B", X"29F", X"2A3", X"2A7", X"2AC", X"2B0", X"2B4", X"2B8", 
X"2BC", X"2C1", X"2C5", X"2C9", X"2CD", X"2D1", X"2D6", X"2DA", X"2DE", X"2E2", 
X"2E6", X"2EA", X"2EF", X"2F3", X"2F7", X"2FB", X"2FF", X"303", X"307", X"30C", 
X"310", X"314", X"318", X"31C", X"320", X"324", X"328", X"32D", X"331", X"335", 
X"339", X"33D", X"341", X"345", X"349", X"34D", X"351", X"355", X"359", X"35D", 
X"362", X"366", X"36A", X"36E", X"372", X"376", X"37A", X"37E", X"382", X"386", 
X"38A", X"38E", X"392", X"396", X"39A", X"39E", X"3A2", X"3A6", X"3AA", X"3AE", 
X"3B2", X"3B6", X"3BA", X"3BE", X"3C1", X"3C5", X"3C9", X"3CD", X"3D1", X"3D5", 
X"3D9", X"3DD", X"3E1", X"3E5", X"3E9", X"3ED", X"3F0", X"3F4", X"3F8", X"3FC", 
X"400", X"404", X"408", X"40C", X"40F", X"413", X"417", X"41B", X"41F", X"423", 
X"426", X"42A", X"42E", X"432", X"436", X"439", X"43D", X"441", X"445", X"449", 
X"44C", X"450", X"454", X"458", X"45B", X"45F", X"463", X"467", X"46A", X"46E", 
X"472", X"476", X"479", X"47D", X"481", X"484", X"488", X"48C", X"48F", X"493", 
X"497", X"49A", X"49E", X"4A2", X"4A5", X"4A9", X"4AD", X"4B0", X"4B4", X"4B7", 
X"4BB", X"4BF", X"4C2", X"4C6", X"4C9", X"4CD", X"4D1", X"4D4", X"4D8", X"4DB", 
X"4DF", X"4E2", X"4E6", X"4E9", X"4ED", X"4F0", X"4F4", X"4F7", X"4FB", X"4FE", 
X"502", X"505", X"509", X"50C", X"510", X"513", X"517", X"51A", X"51E", X"521", 
X"524", X"528", X"52B", X"52F", X"532", X"535", X"539", X"53C", X"540", X"543", 
X"546", X"54A", X"54D", X"550", X"554", X"557", X"55A", X"55E", X"561", X"564", 
X"568", X"56B", X"56E", X"571", X"575", X"578", X"57B", X"57F", X"582", X"585", 
X"588", X"58B", X"58F", X"592", X"595", X"598", X"59B", X"59F", X"5A2", X"5A5", 
X"5A8", X"5AB", X"5AE", X"5B2", X"5B5", X"5B8", X"5BB", X"5BE", X"5C1", X"5C4", 
X"5C7", X"5CA", X"5CE", X"5D1", X"5D4", X"5D7", X"5DA", X"5DD", X"5E0", X"5E3", 
X"5E6", X"5E9", X"5EC", X"5EF", X"5F2", X"5F5", X"5F8", X"5FB", X"5FE", X"601", 
X"604", X"607", X"60A", X"60D", X"60F", X"612", X"615", X"618", X"61B", X"61E", 
X"621", X"624", X"627", X"629", X"62C", X"62F", X"632", X"635", X"638", X"63A", 
X"63D", X"640", X"643", X"646", X"648", X"64B", X"64E", X"651", X"653", X"656", 
X"659", X"65C", X"65E", X"661", X"664", X"666", X"669", X"66C", X"66E", X"671", 
X"674", X"676", X"679", X"67B", X"67E", X"681", X"683", X"686", X"688", X"68B", 
X"68E", X"690", X"693", X"695", X"698", X"69A", X"69D", X"69F", X"6A2", X"6A4", 
X"6A7", X"6A9", X"6AC", X"6AE", X"6B1", X"6B3", X"6B6", X"6B8", X"6BA", X"6BD", 
X"6BF", X"6C2", X"6C4", X"6C6", X"6C9", X"6CB", X"6CE", X"6D0", X"6D2", X"6D5", 
X"6D7", X"6D9", X"6DB", X"6DE", X"6E0", X"6E2", X"6E5", X"6E7", X"6E9", X"6EB", 
X"6EE", X"6F0", X"6F2", X"6F4", X"6F6", X"6F9", X"6FB", X"6FD", X"6FF", X"701", 
X"704", X"706", X"708", X"70A", X"70C", X"70E", X"710", X"712", X"714", X"717", 
X"719", X"71B", X"71D", X"71F", X"721", X"723", X"725", X"727", X"729", X"72B", 
X"72D", X"72F", X"731", X"733", X"735", X"737", X"738", X"73A", X"73C", X"73E", 
X"740", X"742", X"744", X"746", X"748", X"749", X"74B", X"74D", X"74F", X"751", 
X"753", X"754", X"756", X"758", X"75A", X"75B", X"75D", X"75F", X"761", X"762", 
X"764", X"766", X"768", X"769", X"76B", X"76D", X"76E", X"770", X"771", X"773", 
X"775", X"776", X"778", X"77A", X"77B", X"77D", X"77E", X"780", X"781", X"783", 
X"784", X"786", X"788", X"789", X"78B", X"78C", X"78D", X"78F", X"790", X"792", 
X"793", X"795", X"796", X"798", X"799", X"79A", X"79C", X"79D", X"79F", X"7A0", 
X"7A1", X"7A3", X"7A4", X"7A5", X"7A7", X"7A8", X"7A9", X"7AA", X"7AC", X"7AD", 
X"7AE", X"7AF", X"7B1", X"7B2", X"7B3", X"7B4", X"7B6", X"7B7", X"7B8", X"7B9", 
X"7BA", X"7BB", X"7BD", X"7BE", X"7BF", X"7C0", X"7C1", X"7C2", X"7C3", X"7C4", 
X"7C5", X"7C6", X"7C7", X"7C8", X"7C9", X"7CB", X"7CC", X"7CD", X"7CE", X"7CE", 
X"7CF", X"7D0", X"7D1", X"7D2", X"7D3", X"7D4", X"7D5", X"7D6", X"7D7", X"7D8", 
X"7D9", X"7DA", X"7DA", X"7DB", X"7DC", X"7DD", X"7DE", X"7DF", X"7DF", X"7E0", 
X"7E1", X"7E2", X"7E2", X"7E3", X"7E4", X"7E5", X"7E5", X"7E6", X"7E7", X"7E7", 
X"7E8", X"7E9", X"7EA", X"7EA", X"7EB", X"7EB", X"7EC", X"7ED", X"7ED", X"7EE", 
X"7EE", X"7EF", X"7F0", X"7F0", X"7F1", X"7F1", X"7F2", X"7F2", X"7F3", X"7F3", 
X"7F4", X"7F4", X"7F5", X"7F5", X"7F6", X"7F6", X"7F7", X"7F7", X"7F7", X"7F8", 
X"7F8", X"7F9", X"7F9", X"7F9", X"7FA", X"7FA", X"7FA", X"7FB", X"7FB", X"7FB", 
X"7FC", X"7FC", X"7FC", X"7FC", X"7FD", X"7FD", X"7FD", X"7FD", X"7FE", X"7FE", 
X"7FE", X"7FE", X"7FE", X"7FF", X"7FF", X"7FF", X"7FF", X"7FF", X"7FF", X"7FF", 
X"800", X"800", X"800", X"800", X"800", X"800", X"800", X"800", X"800", X"800"
);
begin
	process(H)
	begin
		if(H'event and H='1')then
			SINUS <= "0000"&TABLE(TO_INTEGER(UNSIGNED(ANGLE(15 downto 4))));
			COSINUS <= "0000"&TABLE(TO_INTEGER(UNSIGNED(ANGLE(15 downto 4)))+90*8);
		end if;
	end process;
end architecture;