--   _______    __    ______     ______     _____    ________
--  |   ____|  |  |  |   _  \   |   _  \   / __  \  |___  ___|
--  |  |____   |  |  |  |_|  |  |  |_| /  | |  | |     |  |
--  |   ____|  |  |  |       |  |   _  \  | |  | |     |  |
--  |  |____   |  |  |  |\  \   |  |_| |  | |__| |     |  |
--  |_______|  |__|  |__| \__\  |______/   \_____/     |__|
--
-- Module: TABLE_COSINUS
-- But: Infere une ROM avec COSINUS
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity TABLE_COSINUS is Port ( 
	H       : in  STD_LOGIC;
	ANGLE   : in  STD_LOGIC_VECTOR(14 downto 0);
	COSINUS : out STD_LOGIC_VECTOR(15 downto 0)
);
end TABLE_COSINUS;

architecture Behavioral of TABLE_COSINUS is
TYPE tableSinus is array(0 to (360*64-1)) of STD_LOGIC_VECTOR(15 downto 0);
SIGNAL TABLE : tableSinus := (
X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", 
X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", 
X"8000", X"7FFF", X"7FFF", X"7FFF", X"7FFF", X"7FFF", X"7FFF", X"7FFF", X"7FFF", X"7FFF", 
X"7FFF", X"7FFF", X"7FFF", X"7FFF", X"7FFF", X"7FFF", X"7FFE", X"7FFE", X"7FFE", X"7FFE", 
X"7FFE", X"7FFE", X"7FFE", X"7FFE", X"7FFE", X"7FFE", X"7FFD", X"7FFD", X"7FFD", X"7FFD", 
X"7FFD", X"7FFD", X"7FFD", X"7FFD", X"7FFC", X"7FFC", X"7FFC", X"7FFC", X"7FFC", X"7FFC", 
X"7FFC", X"7FFB", X"7FFB", X"7FFB", X"7FFB", X"7FFB", X"7FFB", X"7FFB", X"7FFA", X"7FFA", 
X"7FFA", X"7FFA", X"7FFA", X"7FFA", X"7FF9", X"7FF9", X"7FF9", X"7FF9", X"7FF9", X"7FF8", 
X"7FF8", X"7FF8", X"7FF8", X"7FF8", X"7FF7", X"7FF7", X"7FF7", X"7FF7", X"7FF7", X"7FF6", 
X"7FF6", X"7FF6", X"7FF6", X"7FF5", X"7FF5", X"7FF5", X"7FF5", X"7FF5", X"7FF4", X"7FF4", 
X"7FF4", X"7FF4", X"7FF3", X"7FF3", X"7FF3", X"7FF3", X"7FF2", X"7FF2", X"7FF2", X"7FF2", 
X"7FF1", X"7FF1", X"7FF1", X"7FF0", X"7FF0", X"7FF0", X"7FF0", X"7FEF", X"7FEF", X"7FEF", 
X"7FEE", X"7FEE", X"7FEE", X"7FEE", X"7FED", X"7FED", X"7FED", X"7FEC", X"7FEC", X"7FEC", 
X"7FEB", X"7FEB", X"7FEB", X"7FEA", X"7FEA", X"7FEA", X"7FE9", X"7FE9", X"7FE9", X"7FE8", 
X"7FE8", X"7FE8", X"7FE7", X"7FE7", X"7FE7", X"7FE6", X"7FE6", X"7FE6", X"7FE5", X"7FE5", 
X"7FE5", X"7FE4", X"7FE4", X"7FE3", X"7FE3", X"7FE3", X"7FE2", X"7FE2", X"7FE2", X"7FE1", 
X"7FE1", X"7FE0", X"7FE0", X"7FE0", X"7FDF", X"7FDF", X"7FDE", X"7FDE", X"7FDE", X"7FDD", 
X"7FDD", X"7FDC", X"7FDC", X"7FDC", X"7FDB", X"7FDB", X"7FDA", X"7FDA", X"7FD9", X"7FD9", 
X"7FD9", X"7FD8", X"7FD8", X"7FD7", X"7FD7", X"7FD6", X"7FD6", X"7FD5", X"7FD5", X"7FD4", 
X"7FD4", X"7FD4", X"7FD3", X"7FD3", X"7FD2", X"7FD2", X"7FD1", X"7FD1", X"7FD0", X"7FD0", 
X"7FCF", X"7FCF", X"7FCE", X"7FCE", X"7FCD", X"7FCD", X"7FCC", X"7FCC", X"7FCB", X"7FCB", 
X"7FCA", X"7FCA", X"7FC9", X"7FC9", X"7FC8", X"7FC8", X"7FC7", X"7FC7", X"7FC6", X"7FC6", 
X"7FC5", X"7FC5", X"7FC4", X"7FC3", X"7FC3", X"7FC2", X"7FC2", X"7FC1", X"7FC1", X"7FC0", 
X"7FC0", X"7FBF", X"7FBE", X"7FBE", X"7FBD", X"7FBD", X"7FBC", X"7FBC", X"7FBB", X"7FBA", 
X"7FBA", X"7FB9", X"7FB9", X"7FB8", X"7FB7", X"7FB7", X"7FB6", X"7FB6", X"7FB5", X"7FB4", 
X"7FB4", X"7FB3", X"7FB3", X"7FB2", X"7FB1", X"7FB1", X"7FB0", X"7FB0", X"7FAF", X"7FAE", 
X"7FAE", X"7FAD", X"7FAC", X"7FAC", X"7FAB", X"7FAA", X"7FAA", X"7FA9", X"7FA9", X"7FA8", 
X"7FA7", X"7FA7", X"7FA6", X"7FA5", X"7FA5", X"7FA4", X"7FA3", X"7FA3", X"7FA2", X"7FA1", 
X"7FA1", X"7FA0", X"7F9F", X"7F9E", X"7F9E", X"7F9D", X"7F9C", X"7F9C", X"7F9B", X"7F9A", 
X"7F9A", X"7F99", X"7F98", X"7F97", X"7F97", X"7F96", X"7F95", X"7F95", X"7F94", X"7F93", 
X"7F92", X"7F92", X"7F91", X"7F90", X"7F8F", X"7F8F", X"7F8E", X"7F8D", X"7F8C", X"7F8C", 
X"7F8B", X"7F8A", X"7F89", X"7F89", X"7F88", X"7F87", X"7F86", X"7F86", X"7F85", X"7F84", 
X"7F83", X"7F83", X"7F82", X"7F81", X"7F80", X"7F7F", X"7F7F", X"7F7E", X"7F7D", X"7F7C", 
X"7F7B", X"7F7B", X"7F7A", X"7F79", X"7F78", X"7F77", X"7F77", X"7F76", X"7F75", X"7F74", 
X"7F73", X"7F72", X"7F72", X"7F71", X"7F70", X"7F6F", X"7F6E", X"7F6D", X"7F6D", X"7F6C", 
X"7F6B", X"7F6A", X"7F69", X"7F68", X"7F67", X"7F67", X"7F66", X"7F65", X"7F64", X"7F63", 
X"7F62", X"7F61", X"7F60", X"7F60", X"7F5F", X"7F5E", X"7F5D", X"7F5C", X"7F5B", X"7F5A", 
X"7F59", X"7F58", X"7F58", X"7F57", X"7F56", X"7F55", X"7F54", X"7F53", X"7F52", X"7F51", 
X"7F50", X"7F4F", X"7F4E", X"7F4D", X"7F4C", X"7F4C", X"7F4B", X"7F4A", X"7F49", X"7F48", 
X"7F47", X"7F46", X"7F45", X"7F44", X"7F43", X"7F42", X"7F41", X"7F40", X"7F3F", X"7F3E", 
X"7F3D", X"7F3C", X"7F3B", X"7F3A", X"7F39", X"7F38", X"7F37", X"7F36", X"7F35", X"7F34", 
X"7F33", X"7F32", X"7F31", X"7F30", X"7F2F", X"7F2E", X"7F2D", X"7F2C", X"7F2B", X"7F2A", 
X"7F29", X"7F28", X"7F27", X"7F26", X"7F25", X"7F24", X"7F23", X"7F22", X"7F21", X"7F20", 
X"7F1F", X"7F1E", X"7F1D", X"7F1C", X"7F1B", X"7F1A", X"7F19", X"7F18", X"7F17", X"7F15", 
X"7F14", X"7F13", X"7F12", X"7F11", X"7F10", X"7F0F", X"7F0E", X"7F0D", X"7F0C", X"7F0B", 
X"7F0A", X"7F08", X"7F07", X"7F06", X"7F05", X"7F04", X"7F03", X"7F02", X"7F01", X"7F00", 
X"7EFF", X"7EFD", X"7EFC", X"7EFB", X"7EFA", X"7EF9", X"7EF8", X"7EF7", X"7EF5", X"7EF4", 
X"7EF3", X"7EF2", X"7EF1", X"7EF0", X"7EEF", X"7EED", X"7EEC", X"7EEB", X"7EEA", X"7EE9", 
X"7EE8", X"7EE6", X"7EE5", X"7EE4", X"7EE3", X"7EE2", X"7EE1", X"7EDF", X"7EDE", X"7EDD", 
X"7EDC", X"7EDB", X"7ED9", X"7ED8", X"7ED7", X"7ED6", X"7ED5", X"7ED3", X"7ED2", X"7ED1", 
X"7ED0", X"7ECF", X"7ECD", X"7ECC", X"7ECB", X"7ECA", X"7EC9", X"7EC7", X"7EC6", X"7EC5", 
X"7EC4", X"7EC2", X"7EC1", X"7EC0", X"7EBF", X"7EBD", X"7EBC", X"7EBB", X"7EBA", X"7EB8", 
X"7EB7", X"7EB6", X"7EB5", X"7EB3", X"7EB2", X"7EB1", X"7EAF", X"7EAE", X"7EAD", X"7EAC", 
X"7EAA", X"7EA9", X"7EA8", X"7EA6", X"7EA5", X"7EA4", X"7EA3", X"7EA1", X"7EA0", X"7E9F", 
X"7E9D", X"7E9C", X"7E9B", X"7E99", X"7E98", X"7E97", X"7E95", X"7E94", X"7E93", X"7E91", 
X"7E90", X"7E8F", X"7E8D", X"7E8C", X"7E8B", X"7E89", X"7E88", X"7E87", X"7E85", X"7E84", 
X"7E83", X"7E81", X"7E80", X"7E7F", X"7E7D", X"7E7C", X"7E7A", X"7E79", X"7E78", X"7E76", 
X"7E75", X"7E74", X"7E72", X"7E71", X"7E6F", X"7E6E", X"7E6D", X"7E6B", X"7E6A", X"7E68", 
X"7E67", X"7E66", X"7E64", X"7E63", X"7E61", X"7E60", X"7E5E", X"7E5D", X"7E5C", X"7E5A", 
X"7E59", X"7E57", X"7E56", X"7E54", X"7E53", X"7E52", X"7E50", X"7E4F", X"7E4D", X"7E4C", 
X"7E4A", X"7E49", X"7E47", X"7E46", X"7E44", X"7E43", X"7E42", X"7E40", X"7E3F", X"7E3D", 
X"7E3C", X"7E3A", X"7E39", X"7E37", X"7E36", X"7E34", X"7E33", X"7E31", X"7E30", X"7E2E", 
X"7E2D", X"7E2B", X"7E2A", X"7E28", X"7E27", X"7E25", X"7E24", X"7E22", X"7E21", X"7E1F", 
X"7E1E", X"7E1C", X"7E1B", X"7E19", X"7E17", X"7E16", X"7E14", X"7E13", X"7E11", X"7E10", 
X"7E0E", X"7E0D", X"7E0B", X"7E0A", X"7E08", X"7E06", X"7E05", X"7E03", X"7E02", X"7E00", 
X"7DFF", X"7DFD", X"7DFB", X"7DFA", X"7DF8", X"7DF7", X"7DF5", X"7DF3", X"7DF2", X"7DF0", 
X"7DEF", X"7DED", X"7DEB", X"7DEA", X"7DE8", X"7DE7", X"7DE5", X"7DE3", X"7DE2", X"7DE0", 
X"7DDF", X"7DDD", X"7DDB", X"7DDA", X"7DD8", X"7DD6", X"7DD5", X"7DD3", X"7DD1", X"7DD0", 
X"7DCE", X"7DCD", X"7DCB", X"7DC9", X"7DC8", X"7DC6", X"7DC4", X"7DC3", X"7DC1", X"7DBF", 
X"7DBE", X"7DBC", X"7DBA", X"7DB9", X"7DB7", X"7DB5", X"7DB4", X"7DB2", X"7DB0", X"7DAE", 
X"7DAD", X"7DAB", X"7DA9", X"7DA8", X"7DA6", X"7DA4", X"7DA3", X"7DA1", X"7D9F", X"7D9D", 
X"7D9C", X"7D9A", X"7D98", X"7D97", X"7D95", X"7D93", X"7D91", X"7D90", X"7D8E", X"7D8C", 
X"7D8A", X"7D89", X"7D87", X"7D85", X"7D83", X"7D82", X"7D80", X"7D7E", X"7D7C", X"7D7B", 
X"7D79", X"7D77", X"7D75", X"7D74", X"7D72", X"7D70", X"7D6E", X"7D6C", X"7D6B", X"7D69", 
X"7D67", X"7D65", X"7D63", X"7D62", X"7D60", X"7D5E", X"7D5C", X"7D5A", X"7D59", X"7D57", 
X"7D55", X"7D53", X"7D51", X"7D50", X"7D4E", X"7D4C", X"7D4A", X"7D48", X"7D46", X"7D45", 
X"7D43", X"7D41", X"7D3F", X"7D3D", X"7D3B", X"7D3A", X"7D38", X"7D36", X"7D34", X"7D32", 
X"7D30", X"7D2E", X"7D2C", X"7D2B", X"7D29", X"7D27", X"7D25", X"7D23", X"7D21", X"7D1F", 
X"7D1D", X"7D1C", X"7D1A", X"7D18", X"7D16", X"7D14", X"7D12", X"7D10", X"7D0E", X"7D0C", 
X"7D0A", X"7D09", X"7D07", X"7D05", X"7D03", X"7D01", X"7CFF", X"7CFD", X"7CFB", X"7CF9", 
X"7CF7", X"7CF5", X"7CF3", X"7CF1", X"7CF0", X"7CEE", X"7CEC", X"7CEA", X"7CE8", X"7CE6", 
X"7CE4", X"7CE2", X"7CE0", X"7CDE", X"7CDC", X"7CDA", X"7CD8", X"7CD6", X"7CD4", X"7CD2", 
X"7CD0", X"7CCE", X"7CCC", X"7CCA", X"7CC8", X"7CC6", X"7CC4", X"7CC2", X"7CC0", X"7CBE", 
X"7CBC", X"7CBA", X"7CB8", X"7CB6", X"7CB4", X"7CB2", X"7CB0", X"7CAE", X"7CAC", X"7CAA", 
X"7CA8", X"7CA6", X"7CA4", X"7CA2", X"7CA0", X"7C9E", X"7C9C", X"7C9A", X"7C98", X"7C96", 
X"7C94", X"7C92", X"7C8F", X"7C8D", X"7C8B", X"7C89", X"7C87", X"7C85", X"7C83", X"7C81", 
X"7C7F", X"7C7D", X"7C7B", X"7C79", X"7C77", X"7C75", X"7C72", X"7C70", X"7C6E", X"7C6C", 
X"7C6A", X"7C68", X"7C66", X"7C64", X"7C62", X"7C60", X"7C5D", X"7C5B", X"7C59", X"7C57", 
X"7C55", X"7C53", X"7C51", X"7C4F", X"7C4C", X"7C4A", X"7C48", X"7C46", X"7C44", X"7C42", 
X"7C40", X"7C3D", X"7C3B", X"7C39", X"7C37", X"7C35", X"7C33", X"7C30", X"7C2E", X"7C2C", 
X"7C2A", X"7C28", X"7C26", X"7C23", X"7C21", X"7C1F", X"7C1D", X"7C1B", X"7C19", X"7C16", 
X"7C14", X"7C12", X"7C10", X"7C0E", X"7C0B", X"7C09", X"7C07", X"7C05", X"7C03", X"7C00", 
X"7BFE", X"7BFC", X"7BFA", X"7BF7", X"7BF5", X"7BF3", X"7BF1", X"7BEE", X"7BEC", X"7BEA", 
X"7BE8", X"7BE6", X"7BE3", X"7BE1", X"7BDF", X"7BDD", X"7BDA", X"7BD8", X"7BD6", X"7BD4", 
X"7BD1", X"7BCF", X"7BCD", X"7BCA", X"7BC8", X"7BC6", X"7BC4", X"7BC1", X"7BBF", X"7BBD", 
X"7BBA", X"7BB8", X"7BB6", X"7BB4", X"7BB1", X"7BAF", X"7BAD", X"7BAA", X"7BA8", X"7BA6", 
X"7BA3", X"7BA1", X"7B9F", X"7B9D", X"7B9A", X"7B98", X"7B96", X"7B93", X"7B91", X"7B8F", 
X"7B8C", X"7B8A", X"7B88", X"7B85", X"7B83", X"7B81", X"7B7E", X"7B7C", X"7B79", X"7B77", 
X"7B75", X"7B72", X"7B70", X"7B6E", X"7B6B", X"7B69", X"7B67", X"7B64", X"7B62", X"7B5F", 
X"7B5D", X"7B5B", X"7B58", X"7B56", X"7B53", X"7B51", X"7B4F", X"7B4C", X"7B4A", X"7B47", 
X"7B45", X"7B43", X"7B40", X"7B3E", X"7B3B", X"7B39", X"7B37", X"7B34", X"7B32", X"7B2F", 
X"7B2D", X"7B2A", X"7B28", X"7B26", X"7B23", X"7B21", X"7B1E", X"7B1C", X"7B19", X"7B17", 
X"7B14", X"7B12", X"7B10", X"7B0D", X"7B0B", X"7B08", X"7B06", X"7B03", X"7B01", X"7AFE", 
X"7AFC", X"7AF9", X"7AF7", X"7AF4", X"7AF2", X"7AEF", X"7AED", X"7AEA", X"7AE8", X"7AE5", 
X"7AE3", X"7AE0", X"7ADE", X"7ADB", X"7AD9", X"7AD6", X"7AD4", X"7AD1", X"7ACF", X"7ACC", 
X"7ACA", X"7AC7", X"7AC5", X"7AC2", X"7AC0", X"7ABD", X"7ABB", X"7AB8", X"7AB6", X"7AB3", 
X"7AB0", X"7AAE", X"7AAB", X"7AA9", X"7AA6", X"7AA4", X"7AA1", X"7A9F", X"7A9C", X"7A99", 
X"7A97", X"7A94", X"7A92", X"7A8F", X"7A8D", X"7A8A", X"7A87", X"7A85", X"7A82", X"7A80", 
X"7A7D", X"7A7A", X"7A78", X"7A75", X"7A73", X"7A70", X"7A6D", X"7A6B", X"7A68", X"7A66", 
X"7A63", X"7A60", X"7A5E", X"7A5B", X"7A58", X"7A56", X"7A53", X"7A51", X"7A4E", X"7A4B", 
X"7A49", X"7A46", X"7A43", X"7A41", X"7A3E", X"7A3B", X"7A39", X"7A36", X"7A33", X"7A31", 
X"7A2E", X"7A2B", X"7A29", X"7A26", X"7A23", X"7A21", X"7A1E", X"7A1B", X"7A19", X"7A16", 
X"7A13", X"7A11", X"7A0E", X"7A0B", X"7A09", X"7A06", X"7A03", X"7A01", X"79FE", X"79FB", 
X"79F8", X"79F6", X"79F3", X"79F0", X"79EE", X"79EB", X"79E8", X"79E5", X"79E3", X"79E0", 
X"79DD", X"79DA", X"79D8", X"79D5", X"79D2", X"79CF", X"79CD", X"79CA", X"79C7", X"79C4", 
X"79C2", X"79BF", X"79BC", X"79B9", X"79B7", X"79B4", X"79B1", X"79AE", X"79AC", X"79A9", 
X"79A6", X"79A3", X"79A0", X"799E", X"799B", X"7998", X"7995", X"7993", X"7990", X"798D", 
X"798A", X"7987", X"7985", X"7982", X"797F", X"797C", X"7979", X"7976", X"7974", X"7971", 
X"796E", X"796B", X"7968", X"7966", X"7963", X"7960", X"795D", X"795A", X"7957", X"7954", 
X"7952", X"794F", X"794C", X"7949", X"7946", X"7943", X"7940", X"793E", X"793B", X"7938", 
X"7935", X"7932", X"792F", X"792C", X"7929", X"7927", X"7924", X"7921", X"791E", X"791B", 
X"7918", X"7915", X"7912", X"790F", X"790D", X"790A", X"7907", X"7904", X"7901", X"78FE", 
X"78FB", X"78F8", X"78F5", X"78F2", X"78EF", X"78EC", X"78EA", X"78E7", X"78E4", X"78E1", 
X"78DE", X"78DB", X"78D8", X"78D5", X"78D2", X"78CF", X"78CC", X"78C9", X"78C6", X"78C3", 
X"78C0", X"78BD", X"78BA", X"78B7", X"78B4", X"78B1", X"78AE", X"78AB", X"78A8", X"78A5", 
X"78A3", X"78A0", X"789D", X"789A", X"7897", X"7894", X"7891", X"788E", X"788B", X"7888", 
X"7885", X"7882", X"787E", X"787B", X"7878", X"7875", X"7872", X"786F", X"786C", X"7869", 
X"7866", X"7863", X"7860", X"785D", X"785A", X"7857", X"7854", X"7851", X"784E", X"784B", 
X"7848", X"7845", X"7842", X"783F", X"783C", X"7839", X"7835", X"7832", X"782F", X"782C", 
X"7829", X"7826", X"7823", X"7820", X"781D", X"781A", X"7817", X"7814", X"7810", X"780D", 
X"780A", X"7807", X"7804", X"7801", X"77FE", X"77FB", X"77F8", X"77F4", X"77F1", X"77EE", 
X"77EB", X"77E8", X"77E5", X"77E2", X"77DF", X"77DB", X"77D8", X"77D5", X"77D2", X"77CF", 
X"77CC", X"77C9", X"77C5", X"77C2", X"77BF", X"77BC", X"77B9", X"77B6", X"77B3", X"77AF", 
X"77AC", X"77A9", X"77A6", X"77A3", X"779F", X"779C", X"7799", X"7796", X"7793", X"7790", 
X"778C", X"7789", X"7786", X"7783", X"7780", X"777C", X"7779", X"7776", X"7773", X"7770", 
X"776C", X"7769", X"7766", X"7763", X"775F", X"775C", X"7759", X"7756", X"7753", X"774F", 
X"774C", X"7749", X"7746", X"7742", X"773F", X"773C", X"7739", X"7735", X"7732", X"772F", 
X"772C", X"7728", X"7725", X"7722", X"771E", X"771B", X"7718", X"7715", X"7711", X"770E", 
X"770B", X"7708", X"7704", X"7701", X"76FE", X"76FA", X"76F7", X"76F4", X"76F0", X"76ED", 
X"76EA", X"76E7", X"76E3", X"76E0", X"76DD", X"76D9", X"76D6", X"76D3", X"76CF", X"76CC", 
X"76C9", X"76C5", X"76C2", X"76BF", X"76BB", X"76B8", X"76B5", X"76B1", X"76AE", X"76AB", 
X"76A7", X"76A4", X"76A1", X"769D", X"769A", X"7696", X"7693", X"7690", X"768C", X"7689", 
X"7686", X"7682", X"767F", X"767B", X"7678", X"7675", X"7671", X"766E", X"766B", X"7667", 
X"7664", X"7660", X"765D", X"765A", X"7656", X"7653", X"764F", X"764C", X"7649", X"7645", 
X"7642", X"763E", X"763B", X"7637", X"7634", X"7631", X"762D", X"762A", X"7626", X"7623", 
X"761F", X"761C", X"7618", X"7615", X"7612", X"760E", X"760B", X"7607", X"7604", X"7600", 
X"75FD", X"75F9", X"75F6", X"75F2", X"75EF", X"75EB", X"75E8", X"75E5", X"75E1", X"75DE", 
X"75DA", X"75D7", X"75D3", X"75D0", X"75CC", X"75C9", X"75C5", X"75C2", X"75BE", X"75BB", 
X"75B7", X"75B4", X"75B0", X"75AD", X"75A9", X"75A6", X"75A2", X"759E", X"759B", X"7597", 
X"7594", X"7590", X"758D", X"7589", X"7586", X"7582", X"757F", X"757B", X"7578", X"7574", 
X"7570", X"756D", X"7569", X"7566", X"7562", X"755F", X"755B", X"7558", X"7554", X"7550", 
X"754D", X"7549", X"7546", X"7542", X"753E", X"753B", X"7537", X"7534", X"7530", X"752D", 
X"7529", X"7525", X"7522", X"751E", X"751B", X"7517", X"7513", X"7510", X"750C", X"7508", 
X"7505", X"7501", X"74FE", X"74FA", X"74F6", X"74F3", X"74EF", X"74EB", X"74E8", X"74E4", 
X"74E1", X"74DD", X"74D9", X"74D6", X"74D2", X"74CE", X"74CB", X"74C7", X"74C3", X"74C0", 
X"74BC", X"74B8", X"74B5", X"74B1", X"74AD", X"74AA", X"74A6", X"74A2", X"749F", X"749B", 
X"7497", X"7493", X"7490", X"748C", X"7488", X"7485", X"7481", X"747D", X"747A", X"7476", 
X"7472", X"746E", X"746B", X"7467", X"7463", X"7460", X"745C", X"7458", X"7454", X"7451", 
X"744D", X"7449", X"7446", X"7442", X"743E", X"743A", X"7437", X"7433", X"742F", X"742B", 
X"7428", X"7424", X"7420", X"741C", X"7419", X"7415", X"7411", X"740D", X"7409", X"7406", 
X"7402", X"73FE", X"73FA", X"73F7", X"73F3", X"73EF", X"73EB", X"73E7", X"73E4", X"73E0", 
X"73DC", X"73D8", X"73D4", X"73D1", X"73CD", X"73C9", X"73C5", X"73C1", X"73BE", X"73BA", 
X"73B6", X"73B2", X"73AE", X"73AA", X"73A7", X"73A3", X"739F", X"739B", X"7397", X"7393", 
X"7390", X"738C", X"7388", X"7384", X"7380", X"737C", X"7379", X"7375", X"7371", X"736D", 
X"7369", X"7365", X"7361", X"735D", X"735A", X"7356", X"7352", X"734E", X"734A", X"7346", 
X"7342", X"733E", X"733B", X"7337", X"7333", X"732F", X"732B", X"7327", X"7323", X"731F", 
X"731B", X"7317", X"7314", X"7310", X"730C", X"7308", X"7304", X"7300", X"72FC", X"72F8", 
X"72F4", X"72F0", X"72EC", X"72E8", X"72E4", X"72E0", X"72DD", X"72D9", X"72D5", X"72D1", 
X"72CD", X"72C9", X"72C5", X"72C1", X"72BD", X"72B9", X"72B5", X"72B1", X"72AD", X"72A9", 
X"72A5", X"72A1", X"729D", X"7299", X"7295", X"7291", X"728D", X"7289", X"7285", X"7281", 
X"727D", X"7279", X"7275", X"7271", X"726D", X"7269", X"7265", X"7261", X"725D", X"7259", 
X"7255", X"7251", X"724D", X"7249", X"7245", X"7241", X"723D", X"7239", X"7235", X"7231", 
X"722D", X"7229", X"7225", X"7221", X"721D", X"7219", X"7215", X"7211", X"720D", X"7208", 
X"7204", X"7200", X"71FC", X"71F8", X"71F4", X"71F0", X"71EC", X"71E8", X"71E4", X"71E0", 
X"71DC", X"71D8", X"71D3", X"71CF", X"71CB", X"71C7", X"71C3", X"71BF", X"71BB", X"71B7", 
X"71B3", X"71AF", X"71AB", X"71A6", X"71A2", X"719E", X"719A", X"7196", X"7192", X"718E", 
X"718A", X"7185", X"7181", X"717D", X"7179", X"7175", X"7171", X"716D", X"7168", X"7164", 
X"7160", X"715C", X"7158", X"7154", X"7150", X"714B", X"7147", X"7143", X"713F", X"713B", 
X"7137", X"7132", X"712E", X"712A", X"7126", X"7122", X"711E", X"7119", X"7115", X"7111", 
X"710D", X"7109", X"7104", X"7100", X"70FC", X"70F8", X"70F4", X"70EF", X"70EB", X"70E7", 
X"70E3", X"70DF", X"70DA", X"70D6", X"70D2", X"70CE", X"70C9", X"70C5", X"70C1", X"70BD", 
X"70B9", X"70B4", X"70B0", X"70AC", X"70A8", X"70A3", X"709F", X"709B", X"7097", X"7092", 
X"708E", X"708A", X"7086", X"7081", X"707D", X"7079", X"7075", X"7070", X"706C", X"7068", 
X"7063", X"705F", X"705B", X"7057", X"7052", X"704E", X"704A", X"7045", X"7041", X"703D", 
X"7039", X"7034", X"7030", X"702C", X"7027", X"7023", X"701F", X"701A", X"7016", X"7012", 
X"700D", X"7009", X"7005", X"7001", X"6FFC", X"6FF8", X"6FF4", X"6FEF", X"6FEB", X"6FE7", 
X"6FE2", X"6FDE", X"6FDA", X"6FD5", X"6FD1", X"6FCC", X"6FC8", X"6FC4", X"6FBF", X"6FBB", 
X"6FB7", X"6FB2", X"6FAE", X"6FAA", X"6FA5", X"6FA1", X"6F9C", X"6F98", X"6F94", X"6F8F", 
X"6F8B", X"6F87", X"6F82", X"6F7E", X"6F79", X"6F75", X"6F71", X"6F6C", X"6F68", X"6F63", 
X"6F5F", X"6F5B", X"6F56", X"6F52", X"6F4D", X"6F49", X"6F45", X"6F40", X"6F3C", X"6F37", 
X"6F33", X"6F2E", X"6F2A", X"6F26", X"6F21", X"6F1D", X"6F18", X"6F14", X"6F0F", X"6F0B", 
X"6F06", X"6F02", X"6EFE", X"6EF9", X"6EF5", X"6EF0", X"6EEC", X"6EE7", X"6EE3", X"6EDE", 
X"6EDA", X"6ED5", X"6ED1", X"6ECD", X"6EC8", X"6EC4", X"6EBF", X"6EBB", X"6EB6", X"6EB2", 
X"6EAD", X"6EA9", X"6EA4", X"6EA0", X"6E9B", X"6E97", X"6E92", X"6E8E", X"6E89", X"6E85", 
X"6E80", X"6E7C", X"6E77", X"6E73", X"6E6E", X"6E6A", X"6E65", X"6E61", X"6E5C", X"6E57", 
X"6E53", X"6E4E", X"6E4A", X"6E45", X"6E41", X"6E3C", X"6E38", X"6E33", X"6E2F", X"6E2A", 
X"6E26", X"6E21", X"6E1C", X"6E18", X"6E13", X"6E0F", X"6E0A", X"6E06", X"6E01", X"6DFC", 
X"6DF8", X"6DF3", X"6DEF", X"6DEA", X"6DE6", X"6DE1", X"6DDC", X"6DD8", X"6DD3", X"6DCF", 
X"6DCA", X"6DC5", X"6DC1", X"6DBC", X"6DB8", X"6DB3", X"6DAE", X"6DAA", X"6DA5", X"6DA1", 
X"6D9C", X"6D97", X"6D93", X"6D8E", X"6D8A", X"6D85", X"6D80", X"6D7C", X"6D77", X"6D72", 
X"6D6E", X"6D69", X"6D64", X"6D60", X"6D5B", X"6D57", X"6D52", X"6D4D", X"6D49", X"6D44", 
X"6D3F", X"6D3B", X"6D36", X"6D31", X"6D2D", X"6D28", X"6D23", X"6D1F", X"6D1A", X"6D15", 
X"6D11", X"6D0C", X"6D07", X"6D03", X"6CFE", X"6CF9", X"6CF5", X"6CF0", X"6CEB", X"6CE6", 
X"6CE2", X"6CDD", X"6CD8", X"6CD4", X"6CCF", X"6CCA", X"6CC6", X"6CC1", X"6CBC", X"6CB7", 
X"6CB3", X"6CAE", X"6CA9", X"6CA4", X"6CA0", X"6C9B", X"6C96", X"6C92", X"6C8D", X"6C88", 
X"6C83", X"6C7F", X"6C7A", X"6C75", X"6C70", X"6C6C", X"6C67", X"6C62", X"6C5D", X"6C59", 
X"6C54", X"6C4F", X"6C4A", X"6C46", X"6C41", X"6C3C", X"6C37", X"6C32", X"6C2E", X"6C29", 
X"6C24", X"6C1F", X"6C1B", X"6C16", X"6C11", X"6C0C", X"6C07", X"6C03", X"6BFE", X"6BF9", 
X"6BF4", X"6BEF", X"6BEB", X"6BE6", X"6BE1", X"6BDC", X"6BD7", X"6BD3", X"6BCE", X"6BC9", 
X"6BC4", X"6BBF", X"6BBA", X"6BB6", X"6BB1", X"6BAC", X"6BA7", X"6BA2", X"6B9D", X"6B99", 
X"6B94", X"6B8F", X"6B8A", X"6B85", X"6B80", X"6B7C", X"6B77", X"6B72", X"6B6D", X"6B68", 
X"6B63", X"6B5E", X"6B5A", X"6B55", X"6B50", X"6B4B", X"6B46", X"6B41", X"6B3C", X"6B37", 
X"6B33", X"6B2E", X"6B29", X"6B24", X"6B1F", X"6B1A", X"6B15", X"6B10", X"6B0B", X"6B07", 
X"6B02", X"6AFD", X"6AF8", X"6AF3", X"6AEE", X"6AE9", X"6AE4", X"6ADF", X"6ADA", X"6AD5", 
X"6AD0", X"6ACC", X"6AC7", X"6AC2", X"6ABD", X"6AB8", X"6AB3", X"6AAE", X"6AA9", X"6AA4", 
X"6A9F", X"6A9A", X"6A95", X"6A90", X"6A8B", X"6A86", X"6A81", X"6A7C", X"6A78", X"6A73", 
X"6A6E", X"6A69", X"6A64", X"6A5F", X"6A5A", X"6A55", X"6A50", X"6A4B", X"6A46", X"6A41", 
X"6A3C", X"6A37", X"6A32", X"6A2D", X"6A28", X"6A23", X"6A1E", X"6A19", X"6A14", X"6A0F", 
X"6A0A", X"6A05", X"6A00", X"69FB", X"69F6", X"69F1", X"69EC", X"69E7", X"69E2", X"69DD", 
X"69D8", X"69D3", X"69CE", X"69C9", X"69C4", X"69BF", X"69BA", X"69B5", X"69AF", X"69AA", 
X"69A5", X"69A0", X"699B", X"6996", X"6991", X"698C", X"6987", X"6982", X"697D", X"6978", 
X"6973", X"696E", X"6969", X"6964", X"695F", X"6959", X"6954", X"694F", X"694A", X"6945", 
X"6940", X"693B", X"6936", X"6931", X"692C", X"6927", X"6922", X"691C", X"6917", X"6912", 
X"690D", X"6908", X"6903", X"68FE", X"68F9", X"68F4", X"68EE", X"68E9", X"68E4", X"68DF", 
X"68DA", X"68D5", X"68D0", X"68CB", X"68C5", X"68C0", X"68BB", X"68B6", X"68B1", X"68AC", 
X"68A7", X"68A1", X"689C", X"6897", X"6892", X"688D", X"6888", X"6883", X"687D", X"6878", 
X"6873", X"686E", X"6869", X"6864", X"685E", X"6859", X"6854", X"684F", X"684A", X"6844", 
X"683F", X"683A", X"6835", X"6830", X"682B", X"6825", X"6820", X"681B", X"6816", X"6811", 
X"680B", X"6806", X"6801", X"67FC", X"67F7", X"67F1", X"67EC", X"67E7", X"67E2", X"67DC", 
X"67D7", X"67D2", X"67CD", X"67C8", X"67C2", X"67BD", X"67B8", X"67B3", X"67AD", X"67A8", 
X"67A3", X"679E", X"6798", X"6793", X"678E", X"6789", X"6783", X"677E", X"6779", X"6774", 
X"676E", X"6769", X"6764", X"675F", X"6759", X"6754", X"674F", X"6749", X"6744", X"673F", 
X"673A", X"6734", X"672F", X"672A", X"6724", X"671F", X"671A", X"6715", X"670F", X"670A", 
X"6705", X"66FF", X"66FA", X"66F5", X"66EF", X"66EA", X"66E5", X"66DF", X"66DA", X"66D5", 
X"66D0", X"66CA", X"66C5", X"66C0", X"66BA", X"66B5", X"66B0", X"66AA", X"66A5", X"66A0", 
X"669A", X"6695", X"668F", X"668A", X"6685", X"667F", X"667A", X"6675", X"666F", X"666A", 
X"6665", X"665F", X"665A", X"6655", X"664F", X"664A", X"6644", X"663F", X"663A", X"6634", 
X"662F", X"662A", X"6624", X"661F", X"6619", X"6614", X"660F", X"6609", X"6604", X"65FE", 
X"65F9", X"65F4", X"65EE", X"65E9", X"65E3", X"65DE", X"65D9", X"65D3", X"65CE", X"65C8", 
X"65C3", X"65BD", X"65B8", X"65B3", X"65AD", X"65A8", X"65A2", X"659D", X"6597", X"6592", 
X"658D", X"6587", X"6582", X"657C", X"6577", X"6571", X"656C", X"6566", X"6561", X"655C", 
X"6556", X"6551", X"654B", X"6546", X"6540", X"653B", X"6535", X"6530", X"652A", X"6525", 
X"651F", X"651A", X"6514", X"650F", X"6509", X"6504", X"64FF", X"64F9", X"64F4", X"64EE", 
X"64E9", X"64E3", X"64DE", X"64D8", X"64D3", X"64CD", X"64C8", X"64C2", X"64BC", X"64B7", 
X"64B1", X"64AC", X"64A6", X"64A1", X"649B", X"6496", X"6490", X"648B", X"6485", X"6480", 
X"647A", X"6475", X"646F", X"646A", X"6464", X"645E", X"6459", X"6453", X"644E", X"6448", 
X"6443", X"643D", X"6438", X"6432", X"642D", X"6427", X"6421", X"641C", X"6416", X"6411", 
X"640B", X"6406", X"6400", X"63FA", X"63F5", X"63EF", X"63EA", X"63E4", X"63DE", X"63D9", 
X"63D3", X"63CE", X"63C8", X"63C2", X"63BD", X"63B7", X"63B2", X"63AC", X"63A6", X"63A1", 
X"639B", X"6396", X"6390", X"638A", X"6385", X"637F", X"637A", X"6374", X"636E", X"6369", 
X"6363", X"635D", X"6358", X"6352", X"634C", X"6347", X"6341", X"633C", X"6336", X"6330", 
X"632B", X"6325", X"631F", X"631A", X"6314", X"630E", X"6309", X"6303", X"62FD", X"62F8", 
X"62F2", X"62EC", X"62E7", X"62E1", X"62DB", X"62D6", X"62D0", X"62CA", X"62C5", X"62BF", 
X"62B9", X"62B4", X"62AE", X"62A8", X"62A2", X"629D", X"6297", X"6291", X"628C", X"6286", 
X"6280", X"627B", X"6275", X"626F", X"6269", X"6264", X"625E", X"6258", X"6253", X"624D", 
X"6247", X"6241", X"623C", X"6236", X"6230", X"622A", X"6225", X"621F", X"6219", X"6213", 
X"620E", X"6208", X"6202", X"61FD", X"61F7", X"61F1", X"61EB", X"61E5", X"61E0", X"61DA", 
X"61D4", X"61CE", X"61C9", X"61C3", X"61BD", X"61B7", X"61B2", X"61AC", X"61A6", X"61A0", 
X"619A", X"6195", X"618F", X"6189", X"6183", X"617E", X"6178", X"6172", X"616C", X"6166", 
X"6161", X"615B", X"6155", X"614F", X"6149", X"6144", X"613E", X"6138", X"6132", X"612C", 
X"6126", X"6121", X"611B", X"6115", X"610F", X"6109", X"6104", X"60FE", X"60F8", X"60F2", 
X"60EC", X"60E6", X"60E1", X"60DB", X"60D5", X"60CF", X"60C9", X"60C3", X"60BD", X"60B8", 
X"60B2", X"60AC", X"60A6", X"60A0", X"609A", X"6094", X"608F", X"6089", X"6083", X"607D", 
X"6077", X"6071", X"606B", X"6065", X"6060", X"605A", X"6054", X"604E", X"6048", X"6042", 
X"603C", X"6036", X"6031", X"602B", X"6025", X"601F", X"6019", X"6013", X"600D", X"6007", 
X"6001", X"5FFB", X"5FF5", X"5FF0", X"5FEA", X"5FE4", X"5FDE", X"5FD8", X"5FD2", X"5FCC", 
X"5FC6", X"5FC0", X"5FBA", X"5FB4", X"5FAE", X"5FA8", X"5FA2", X"5F9D", X"5F97", X"5F91", 
X"5F8B", X"5F85", X"5F7F", X"5F79", X"5F73", X"5F6D", X"5F67", X"5F61", X"5F5B", X"5F55", 
X"5F4F", X"5F49", X"5F43", X"5F3D", X"5F37", X"5F31", X"5F2B", X"5F25", X"5F1F", X"5F19", 
X"5F13", X"5F0D", X"5F07", X"5F01", X"5EFB", X"5EF5", X"5EEF", X"5EE9", X"5EE3", X"5EDD", 
X"5ED7", X"5ED1", X"5ECB", X"5EC5", X"5EBF", X"5EB9", X"5EB3", X"5EAD", X"5EA7", X"5EA1", 
X"5E9B", X"5E95", X"5E8F", X"5E89", X"5E83", X"5E7D", X"5E77", X"5E71", X"5E6B", X"5E65", 
X"5E5F", X"5E59", X"5E53", X"5E4D", X"5E47", X"5E41", X"5E3B", X"5E35", X"5E2F", X"5E29", 
X"5E23", X"5E1D", X"5E17", X"5E10", X"5E0A", X"5E04", X"5DFE", X"5DF8", X"5DF2", X"5DEC", 
X"5DE6", X"5DE0", X"5DDA", X"5DD4", X"5DCE", X"5DC8", X"5DC2", X"5DBB", X"5DB5", X"5DAF", 
X"5DA9", X"5DA3", X"5D9D", X"5D97", X"5D91", X"5D8B", X"5D85", X"5D7F", X"5D78", X"5D72", 
X"5D6C", X"5D66", X"5D60", X"5D5A", X"5D54", X"5D4E", X"5D48", X"5D41", X"5D3B", X"5D35", 
X"5D2F", X"5D29", X"5D23", X"5D1D", X"5D16", X"5D10", X"5D0A", X"5D04", X"5CFE", X"5CF8", 
X"5CF2", X"5CEC", X"5CE5", X"5CDF", X"5CD9", X"5CD3", X"5CCD", X"5CC7", X"5CC0", X"5CBA", 
X"5CB4", X"5CAE", X"5CA8", X"5CA2", X"5C9B", X"5C95", X"5C8F", X"5C89", X"5C83", X"5C7D", 
X"5C76", X"5C70", X"5C6A", X"5C64", X"5C5E", X"5C58", X"5C51", X"5C4B", X"5C45", X"5C3F", 
X"5C39", X"5C32", X"5C2C", X"5C26", X"5C20", X"5C1A", X"5C13", X"5C0D", X"5C07", X"5C01", 
X"5BFA", X"5BF4", X"5BEE", X"5BE8", X"5BE2", X"5BDB", X"5BD5", X"5BCF", X"5BC9", X"5BC2", 
X"5BBC", X"5BB6", X"5BB0", X"5BAA", X"5BA3", X"5B9D", X"5B97", X"5B91", X"5B8A", X"5B84", 
X"5B7E", X"5B78", X"5B71", X"5B6B", X"5B65", X"5B5F", X"5B58", X"5B52", X"5B4C", X"5B46", 
X"5B3F", X"5B39", X"5B33", X"5B2C", X"5B26", X"5B20", X"5B1A", X"5B13", X"5B0D", X"5B07", 
X"5B01", X"5AFA", X"5AF4", X"5AEE", X"5AE7", X"5AE1", X"5ADB", X"5AD4", X"5ACE", X"5AC8", 
X"5AC2", X"5ABB", X"5AB5", X"5AAF", X"5AA8", X"5AA2", X"5A9C", X"5A95", X"5A8F", X"5A89", 
X"5A82", X"5A7C", X"5A76", X"5A70", X"5A69", X"5A63", X"5A5D", X"5A56", X"5A50", X"5A4A", 
X"5A43", X"5A3D", X"5A37", X"5A30", X"5A2A", X"5A24", X"5A1D", X"5A17", X"5A10", X"5A0A", 
X"5A04", X"59FD", X"59F7", X"59F1", X"59EA", X"59E4", X"59DE", X"59D7", X"59D1", X"59CB", 
X"59C4", X"59BE", X"59B7", X"59B1", X"59AB", X"59A4", X"599E", X"5998", X"5991", X"598B", 
X"5984", X"597E", X"5978", X"5971", X"596B", X"5964", X"595E", X"5958", X"5951", X"594B", 
X"5944", X"593E", X"5938", X"5931", X"592B", X"5924", X"591E", X"5918", X"5911", X"590B", 
X"5904", X"58FE", X"58F7", X"58F1", X"58EB", X"58E4", X"58DE", X"58D7", X"58D1", X"58CA", 
X"58C4", X"58BE", X"58B7", X"58B1", X"58AA", X"58A4", X"589D", X"5897", X"5890", X"588A", 
X"5884", X"587D", X"5877", X"5870", X"586A", X"5863", X"585D", X"5856", X"5850", X"5849", 
X"5843", X"583C", X"5836", X"582F", X"5829", X"5822", X"581C", X"5816", X"580F", X"5809", 
X"5802", X"57FC", X"57F5", X"57EF", X"57E8", X"57E2", X"57DB", X"57D5", X"57CE", X"57C8", 
X"57C1", X"57BB", X"57B4", X"57AE", X"57A7", X"57A1", X"579A", X"5794", X"578D", X"5786", 
X"5780", X"5779", X"5773", X"576C", X"5766", X"575F", X"5759", X"5752", X"574C", X"5745", 
X"573F", X"5738", X"5732", X"572B", X"5724", X"571E", X"5717", X"5711", X"570A", X"5704", 
X"56FD", X"56F7", X"56F0", X"56EA", X"56E3", X"56DC", X"56D6", X"56CF", X"56C9", X"56C2", 
X"56BC", X"56B5", X"56AE", X"56A8", X"56A1", X"569B", X"5694", X"568D", X"5687", X"5680", 
X"567A", X"5673", X"566D", X"5666", X"565F", X"5659", X"5652", X"564C", X"5645", X"563E", 
X"5638", X"5631", X"562B", X"5624", X"561D", X"5617", X"5610", X"560A", X"5603", X"55FC", 
X"55F6", X"55EF", X"55E8", X"55E2", X"55DB", X"55D5", X"55CE", X"55C7", X"55C1", X"55BA", 
X"55B3", X"55AD", X"55A6", X"559F", X"5599", X"5592", X"558B", X"5585", X"557E", X"5578", 
X"5571", X"556A", X"5564", X"555D", X"5556", X"5550", X"5549", X"5542", X"553C", X"5535", 
X"552E", X"5528", X"5521", X"551A", X"5514", X"550D", X"5506", X"5500", X"54F9", X"54F2", 
X"54EB", X"54E5", X"54DE", X"54D7", X"54D1", X"54CA", X"54C3", X"54BD", X"54B6", X"54AF", 
X"54A9", X"54A2", X"549B", X"5494", X"548E", X"5487", X"5480", X"547A", X"5473", X"546C", 
X"5465", X"545F", X"5458", X"5451", X"544B", X"5444", X"543D", X"5436", X"5430", X"5429", 
X"5422", X"541B", X"5415", X"540E", X"5407", X"5400", X"53FA", X"53F3", X"53EC", X"53E6", 
X"53DF", X"53D8", X"53D1", X"53CA", X"53C4", X"53BD", X"53B6", X"53AF", X"53A9", X"53A2", 
X"539B", X"5394", X"538E", X"5387", X"5380", X"5379", X"5373", X"536C", X"5365", X"535E", 
X"5357", X"5351", X"534A", X"5343", X"533C", X"5335", X"532F", X"5328", X"5321", X"531A", 
X"5314", X"530D", X"5306", X"52FF", X"52F8", X"52F2", X"52EB", X"52E4", X"52DD", X"52D6", 
X"52CF", X"52C9", X"52C2", X"52BB", X"52B4", X"52AD", X"52A7", X"52A0", X"5299", X"5292", 
X"528B", X"5284", X"527E", X"5277", X"5270", X"5269", X"5262", X"525B", X"5255", X"524E", 
X"5247", X"5240", X"5239", X"5232", X"522B", X"5225", X"521E", X"5217", X"5210", X"5209", 
X"5202", X"51FB", X"51F5", X"51EE", X"51E7", X"51E0", X"51D9", X"51D2", X"51CB", X"51C5", 
X"51BE", X"51B7", X"51B0", X"51A9", X"51A2", X"519B", X"5194", X"518D", X"5187", X"5180", 
X"5179", X"5172", X"516B", X"5164", X"515D", X"5156", X"514F", X"5149", X"5142", X"513B", 
X"5134", X"512D", X"5126", X"511F", X"5118", X"5111", X"510A", X"5103", X"50FC", X"50F6", 
X"50EF", X"50E8", X"50E1", X"50DA", X"50D3", X"50CC", X"50C5", X"50BE", X"50B7", X"50B0", 
X"50A9", X"50A2", X"509B", X"5095", X"508E", X"5087", X"5080", X"5079", X"5072", X"506B", 
X"5064", X"505D", X"5056", X"504F", X"5048", X"5041", X"503A", X"5033", X"502C", X"5025", 
X"501E", X"5017", X"5010", X"5009", X"5002", X"4FFB", X"4FF4", X"4FED", X"4FE6", X"4FDF", 
X"4FD8", X"4FD2", X"4FCB", X"4FC4", X"4FBD", X"4FB6", X"4FAF", X"4FA8", X"4FA1", X"4F9A", 
X"4F93", X"4F8C", X"4F85", X"4F7E", X"4F77", X"4F70", X"4F69", X"4F62", X"4F5B", X"4F54", 
X"4F4D", X"4F45", X"4F3E", X"4F37", X"4F30", X"4F29", X"4F22", X"4F1B", X"4F14", X"4F0D", 
X"4F06", X"4EFF", X"4EF8", X"4EF1", X"4EEA", X"4EE3", X"4EDC", X"4ED5", X"4ECE", X"4EC7", 
X"4EC0", X"4EB9", X"4EB2", X"4EAB", X"4EA4", X"4E9D", X"4E96", X"4E8F", X"4E88", X"4E80", 
X"4E79", X"4E72", X"4E6B", X"4E64", X"4E5D", X"4E56", X"4E4F", X"4E48", X"4E41", X"4E3A", 
X"4E33", X"4E2C", X"4E25", X"4E1D", X"4E16", X"4E0F", X"4E08", X"4E01", X"4DFA", X"4DF3", 
X"4DEC", X"4DE5", X"4DDE", X"4DD7", X"4DD0", X"4DC8", X"4DC1", X"4DBA", X"4DB3", X"4DAC", 
X"4DA5", X"4D9E", X"4D97", X"4D90", X"4D88", X"4D81", X"4D7A", X"4D73", X"4D6C", X"4D65", 
X"4D5E", X"4D57", X"4D50", X"4D48", X"4D41", X"4D3A", X"4D33", X"4D2C", X"4D25", X"4D1E", 
X"4D17", X"4D0F", X"4D08", X"4D01", X"4CFA", X"4CF3", X"4CEC", X"4CE5", X"4CDD", X"4CD6", 
X"4CCF", X"4CC8", X"4CC1", X"4CBA", X"4CB3", X"4CAB", X"4CA4", X"4C9D", X"4C96", X"4C8F", 
X"4C88", X"4C80", X"4C79", X"4C72", X"4C6B", X"4C64", X"4C5D", X"4C55", X"4C4E", X"4C47", 
X"4C40", X"4C39", X"4C32", X"4C2A", X"4C23", X"4C1C", X"4C15", X"4C0E", X"4C06", X"4BFF", 
X"4BF8", X"4BF1", X"4BEA", X"4BE2", X"4BDB", X"4BD4", X"4BCD", X"4BC6", X"4BBE", X"4BB7", 
X"4BB0", X"4BA9", X"4BA2", X"4B9A", X"4B93", X"4B8C", X"4B85", X"4B7E", X"4B76", X"4B6F", 
X"4B68", X"4B61", X"4B59", X"4B52", X"4B4B", X"4B44", X"4B3D", X"4B35", X"4B2E", X"4B27", 
X"4B20", X"4B18", X"4B11", X"4B0A", X"4B03", X"4AFB", X"4AF4", X"4AED", X"4AE6", X"4ADE", 
X"4AD7", X"4AD0", X"4AC9", X"4AC1", X"4ABA", X"4AB3", X"4AAC", X"4AA4", X"4A9D", X"4A96", 
X"4A8F", X"4A87", X"4A80", X"4A79", X"4A72", X"4A6A", X"4A63", X"4A5C", X"4A54", X"4A4D", 
X"4A46", X"4A3F", X"4A37", X"4A30", X"4A29", X"4A22", X"4A1A", X"4A13", X"4A0C", X"4A04", 
X"49FD", X"49F6", X"49EE", X"49E7", X"49E0", X"49D9", X"49D1", X"49CA", X"49C3", X"49BB", 
X"49B4", X"49AD", X"49A5", X"499E", X"4997", X"4990", X"4988", X"4981", X"497A", X"4972", 
X"496B", X"4964", X"495C", X"4955", X"494E", X"4946", X"493F", X"4938", X"4930", X"4929", 
X"4922", X"491A", X"4913", X"490C", X"4904", X"48FD", X"48F6", X"48EE", X"48E7", X"48E0", 
X"48D8", X"48D1", X"48CA", X"48C2", X"48BB", X"48B4", X"48AC", X"48A5", X"489D", X"4896", 
X"488F", X"4887", X"4880", X"4879", X"4871", X"486A", X"4863", X"485B", X"4854", X"484C", 
X"4845", X"483E", X"4836", X"482F", X"4828", X"4820", X"4819", X"4811", X"480A", X"4803", 
X"47FB", X"47F4", X"47EC", X"47E5", X"47DE", X"47D6", X"47CF", X"47C7", X"47C0", X"47B9", 
X"47B1", X"47AA", X"47A2", X"479B", X"4794", X"478C", X"4785", X"477D", X"4776", X"476F", 
X"4767", X"4760", X"4758", X"4751", X"4749", X"4742", X"473B", X"4733", X"472C", X"4724", 
X"471D", X"4715", X"470E", X"4707", X"46FF", X"46F8", X"46F0", X"46E9", X"46E1", X"46DA", 
X"46D3", X"46CB", X"46C4", X"46BC", X"46B5", X"46AD", X"46A6", X"469E", X"4697", X"4690", 
X"4688", X"4681", X"4679", X"4672", X"466A", X"4663", X"465B", X"4654", X"464C", X"4645", 
X"463D", X"4636", X"462E", X"4627", X"4620", X"4618", X"4611", X"4609", X"4602", X"45FA", 
X"45F3", X"45EB", X"45E4", X"45DC", X"45D5", X"45CD", X"45C6", X"45BE", X"45B7", X"45AF", 
X"45A8", X"45A0", X"4599", X"4591", X"458A", X"4582", X"457B", X"4573", X"456C", X"4564", 
X"455D", X"4555", X"454E", X"4546", X"453F", X"4537", X"4530", X"4528", X"4521", X"4519", 
X"4512", X"450A", X"4502", X"44FB", X"44F3", X"44EC", X"44E4", X"44DD", X"44D5", X"44CE", 
X"44C6", X"44BF", X"44B7", X"44B0", X"44A8", X"44A1", X"4499", X"4491", X"448A", X"4482", 
X"447B", X"4473", X"446C", X"4464", X"445D", X"4455", X"444D", X"4446", X"443E", X"4437", 
X"442F", X"4428", X"4420", X"4419", X"4411", X"4409", X"4402", X"43FA", X"43F3", X"43EB", 
X"43E4", X"43DC", X"43D4", X"43CD", X"43C5", X"43BE", X"43B6", X"43AE", X"43A7", X"439F", 
X"4398", X"4390", X"4389", X"4381", X"4379", X"4372", X"436A", X"4363", X"435B", X"4353", 
X"434C", X"4344", X"433D", X"4335", X"432D", X"4326", X"431E", X"4317", X"430F", X"4307", 
X"4300", X"42F8", X"42F0", X"42E9", X"42E1", X"42DA", X"42D2", X"42CA", X"42C3", X"42BB", 
X"42B3", X"42AC", X"42A4", X"429D", X"4295", X"428D", X"4286", X"427E", X"4276", X"426F", 
X"4267", X"4260", X"4258", X"4250", X"4249", X"4241", X"4239", X"4232", X"422A", X"4222", 
X"421B", X"4213", X"420B", X"4204", X"41FC", X"41F4", X"41ED", X"41E5", X"41DD", X"41D6", 
X"41CE", X"41C6", X"41BF", X"41B7", X"41AF", X"41A8", X"41A0", X"4198", X"4191", X"4189", 
X"4181", X"417A", X"4172", X"416A", X"4163", X"415B", X"4153", X"414C", X"4144", X"413C", 
X"4135", X"412D", X"4125", X"411E", X"4116", X"410E", X"4106", X"40FF", X"40F7", X"40EF", 
X"40E8", X"40E0", X"40D8", X"40D1", X"40C9", X"40C1", X"40B9", X"40B2", X"40AA", X"40A2", 
X"409B", X"4093", X"408B", X"4083", X"407C", X"4074", X"406C", X"4065", X"405D", X"4055", 
X"404D", X"4046", X"403E", X"4036", X"402E", X"4027", X"401F", X"4017", X"400F", X"4008", 
X"4000", X"3FF8", X"3FF1", X"3FE9", X"3FE1", X"3FD9", X"3FD2", X"3FCA", X"3FC2", X"3FBA", 
X"3FB3", X"3FAB", X"3FA3", X"3F9B", X"3F94", X"3F8C", X"3F84", X"3F7C", X"3F75", X"3F6D", 
X"3F65", X"3F5D", X"3F55", X"3F4E", X"3F46", X"3F3E", X"3F36", X"3F2F", X"3F27", X"3F1F", 
X"3F17", X"3F10", X"3F08", X"3F00", X"3EF8", X"3EF0", X"3EE9", X"3EE1", X"3ED9", X"3ED1", 
X"3EC9", X"3EC2", X"3EBA", X"3EB2", X"3EAA", X"3EA3", X"3E9B", X"3E93", X"3E8B", X"3E83", 
X"3E7C", X"3E74", X"3E6C", X"3E64", X"3E5C", X"3E55", X"3E4D", X"3E45", X"3E3D", X"3E35", 
X"3E2D", X"3E26", X"3E1E", X"3E16", X"3E0E", X"3E06", X"3DFF", X"3DF7", X"3DEF", X"3DE7", 
X"3DDF", X"3DD8", X"3DD0", X"3DC8", X"3DC0", X"3DB8", X"3DB0", X"3DA9", X"3DA1", X"3D99", 
X"3D91", X"3D89", X"3D81", X"3D7A", X"3D72", X"3D6A", X"3D62", X"3D5A", X"3D52", X"3D4A", 
X"3D43", X"3D3B", X"3D33", X"3D2B", X"3D23", X"3D1B", X"3D14", X"3D0C", X"3D04", X"3CFC", 
X"3CF4", X"3CEC", X"3CE4", X"3CDD", X"3CD5", X"3CCD", X"3CC5", X"3CBD", X"3CB5", X"3CAD", 
X"3CA5", X"3C9E", X"3C96", X"3C8E", X"3C86", X"3C7E", X"3C76", X"3C6E", X"3C66", X"3C5F", 
X"3C57", X"3C4F", X"3C47", X"3C3F", X"3C37", X"3C2F", X"3C27", X"3C20", X"3C18", X"3C10", 
X"3C08", X"3C00", X"3BF8", X"3BF0", X"3BE8", X"3BE0", X"3BD8", X"3BD1", X"3BC9", X"3BC1", 
X"3BB9", X"3BB1", X"3BA9", X"3BA1", X"3B99", X"3B91", X"3B89", X"3B82", X"3B7A", X"3B72", 
X"3B6A", X"3B62", X"3B5A", X"3B52", X"3B4A", X"3B42", X"3B3A", X"3B32", X"3B2A", X"3B23", 
X"3B1B", X"3B13", X"3B0B", X"3B03", X"3AFB", X"3AF3", X"3AEB", X"3AE3", X"3ADB", X"3AD3", 
X"3ACB", X"3AC3", X"3ABB", X"3AB3", X"3AAB", X"3AA4", X"3A9C", X"3A94", X"3A8C", X"3A84", 
X"3A7C", X"3A74", X"3A6C", X"3A64", X"3A5C", X"3A54", X"3A4C", X"3A44", X"3A3C", X"3A34", 
X"3A2C", X"3A24", X"3A1C", X"3A14", X"3A0C", X"3A04", X"39FD", X"39F5", X"39ED", X"39E5", 
X"39DD", X"39D5", X"39CD", X"39C5", X"39BD", X"39B5", X"39AD", X"39A5", X"399D", X"3995", 
X"398D", X"3985", X"397D", X"3975", X"396D", X"3965", X"395D", X"3955", X"394D", X"3945", 
X"393D", X"3935", X"392D", X"3925", X"391D", X"3915", X"390D", X"3905", X"38FD", X"38F5", 
X"38ED", X"38E5", X"38DD", X"38D5", X"38CD", X"38C5", X"38BD", X"38B5", X"38AD", X"38A5", 
X"389D", X"3895", X"388D", X"3885", X"387D", X"3875", X"386D", X"3865", X"385D", X"3855", 
X"384D", X"3845", X"383D", X"3835", X"382D", X"3825", X"381D", X"3815", X"380C", X"3804", 
X"37FC", X"37F4", X"37EC", X"37E4", X"37DC", X"37D4", X"37CC", X"37C4", X"37BC", X"37B4", 
X"37AC", X"37A4", X"379C", X"3794", X"378C", X"3784", X"377C", X"3774", X"376C", X"3764", 
X"375B", X"3753", X"374B", X"3743", X"373B", X"3733", X"372B", X"3723", X"371B", X"3713", 
X"370B", X"3703", X"36FB", X"36F3", X"36EB", X"36E3", X"36DA", X"36D2", X"36CA", X"36C2", 
X"36BA", X"36B2", X"36AA", X"36A2", X"369A", X"3692", X"368A", X"3682", X"3679", X"3671", 
X"3669", X"3661", X"3659", X"3651", X"3649", X"3641", X"3639", X"3631", X"3629", X"3620", 
X"3618", X"3610", X"3608", X"3600", X"35F8", X"35F0", X"35E8", X"35E0", X"35D8", X"35CF", 
X"35C7", X"35BF", X"35B7", X"35AF", X"35A7", X"359F", X"3597", X"358F", X"3586", X"357E", 
X"3576", X"356E", X"3566", X"355E", X"3556", X"354E", X"3545", X"353D", X"3535", X"352D", 
X"3525", X"351D", X"3515", X"350D", X"3504", X"34FC", X"34F4", X"34EC", X"34E4", X"34DC", 
X"34D4", X"34CB", X"34C3", X"34BB", X"34B3", X"34AB", X"34A3", X"349B", X"3492", X"348A", 
X"3482", X"347A", X"3472", X"346A", X"3462", X"3459", X"3451", X"3449", X"3441", X"3439", 
X"3431", X"3428", X"3420", X"3418", X"3410", X"3408", X"3400", X"33F7", X"33EF", X"33E7", 
X"33DF", X"33D7", X"33CF", X"33C6", X"33BE", X"33B6", X"33AE", X"33A6", X"339E", X"3395", 
X"338D", X"3385", X"337D", X"3375", X"336C", X"3364", X"335C", X"3354", X"334C", X"3344", 
X"333B", X"3333", X"332B", X"3323", X"331B", X"3312", X"330A", X"3302", X"32FA", X"32F2", 
X"32E9", X"32E1", X"32D9", X"32D1", X"32C9", X"32C0", X"32B8", X"32B0", X"32A8", X"32A0", 
X"3297", X"328F", X"3287", X"327F", X"3277", X"326E", X"3266", X"325E", X"3256", X"324D", 
X"3245", X"323D", X"3235", X"322D", X"3224", X"321C", X"3214", X"320C", X"3203", X"31FB", 
X"31F3", X"31EB", X"31E3", X"31DA", X"31D2", X"31CA", X"31C2", X"31B9", X"31B1", X"31A9", 
X"31A1", X"3198", X"3190", X"3188", X"3180", X"3178", X"316F", X"3167", X"315F", X"3157", 
X"314E", X"3146", X"313E", X"3136", X"312D", X"3125", X"311D", X"3115", X"310C", X"3104", 
X"30FC", X"30F4", X"30EB", X"30E3", X"30DB", X"30D2", X"30CA", X"30C2", X"30BA", X"30B1", 
X"30A9", X"30A1", X"3099", X"3090", X"3088", X"3080", X"3078", X"306F", X"3067", X"305F", 
X"3056", X"304E", X"3046", X"303E", X"3035", X"302D", X"3025", X"301D", X"3014", X"300C", 
X"3004", X"2FFB", X"2FF3", X"2FEB", X"2FE3", X"2FDA", X"2FD2", X"2FCA", X"2FC1", X"2FB9", 
X"2FB1", X"2FA9", X"2FA0", X"2F98", X"2F90", X"2F87", X"2F7F", X"2F77", X"2F6E", X"2F66", 
X"2F5E", X"2F56", X"2F4D", X"2F45", X"2F3D", X"2F34", X"2F2C", X"2F24", X"2F1B", X"2F13", 
X"2F0B", X"2F02", X"2EFA", X"2EF2", X"2EEA", X"2EE1", X"2ED9", X"2ED1", X"2EC8", X"2EC0", 
X"2EB8", X"2EAF", X"2EA7", X"2E9F", X"2E96", X"2E8E", X"2E86", X"2E7D", X"2E75", X"2E6D", 
X"2E64", X"2E5C", X"2E54", X"2E4B", X"2E43", X"2E3B", X"2E32", X"2E2A", X"2E22", X"2E19", 
X"2E11", X"2E09", X"2E00", X"2DF8", X"2DF0", X"2DE7", X"2DDF", X"2DD7", X"2DCE", X"2DC6", 
X"2DBE", X"2DB5", X"2DAD", X"2DA5", X"2D9C", X"2D94", X"2D8C", X"2D83", X"2D7B", X"2D72", 
X"2D6A", X"2D62", X"2D59", X"2D51", X"2D49", X"2D40", X"2D38", X"2D30", X"2D27", X"2D1F", 
X"2D17", X"2D0E", X"2D06", X"2CFD", X"2CF5", X"2CED", X"2CE4", X"2CDC", X"2CD4", X"2CCB", 
X"2CC3", X"2CBA", X"2CB2", X"2CAA", X"2CA1", X"2C99", X"2C91", X"2C88", X"2C80", X"2C77", 
X"2C6F", X"2C67", X"2C5E", X"2C56", X"2C4E", X"2C45", X"2C3D", X"2C34", X"2C2C", X"2C24", 
X"2C1B", X"2C13", X"2C0A", X"2C02", X"2BFA", X"2BF1", X"2BE9", X"2BE1", X"2BD8", X"2BD0", 
X"2BC7", X"2BBF", X"2BB7", X"2BAE", X"2BA6", X"2B9D", X"2B95", X"2B8D", X"2B84", X"2B7C", 
X"2B73", X"2B6B", X"2B62", X"2B5A", X"2B52", X"2B49", X"2B41", X"2B38", X"2B30", X"2B28", 
X"2B1F", X"2B17", X"2B0E", X"2B06", X"2AFE", X"2AF5", X"2AED", X"2AE4", X"2ADC", X"2AD3", 
X"2ACB", X"2AC3", X"2ABA", X"2AB2", X"2AA9", X"2AA1", X"2A98", X"2A90", X"2A88", X"2A7F", 
X"2A77", X"2A6E", X"2A66", X"2A5D", X"2A55", X"2A4D", X"2A44", X"2A3C", X"2A33", X"2A2B", 
X"2A22", X"2A1A", X"2A12", X"2A09", X"2A01", X"29F8", X"29F0", X"29E7", X"29DF", X"29D6", 
X"29CE", X"29C6", X"29BD", X"29B5", X"29AC", X"29A4", X"299B", X"2993", X"298A", X"2982", 
X"297A", X"2971", X"2969", X"2960", X"2958", X"294F", X"2947", X"293E", X"2936", X"292D", 
X"2925", X"291C", X"2914", X"290C", X"2903", X"28FB", X"28F2", X"28EA", X"28E1", X"28D9", 
X"28D0", X"28C8", X"28BF", X"28B7", X"28AE", X"28A6", X"289D", X"2895", X"288C", X"2884", 
X"287C", X"2873", X"286B", X"2862", X"285A", X"2851", X"2849", X"2840", X"2838", X"282F", 
X"2827", X"281E", X"2816", X"280D", X"2805", X"27FC", X"27F4", X"27EB", X"27E3", X"27DA", 
X"27D2", X"27C9", X"27C1", X"27B8", X"27B0", X"27A7", X"279F", X"2796", X"278E", X"2785", 
X"277D", X"2774", X"276C", X"2763", X"275B", X"2752", X"274A", X"2741", X"2739", X"2730", 
X"2728", X"271F", X"2717", X"270E", X"2706", X"26FD", X"26F5", X"26EC", X"26E4", X"26DB", 
X"26D3", X"26CA", X"26C2", X"26B9", X"26B1", X"26A8", X"26A0", X"2697", X"268F", X"2686", 
X"267E", X"2675", X"266C", X"2664", X"265B", X"2653", X"264A", X"2642", X"2639", X"2631", 
X"2628", X"2620", X"2617", X"260F", X"2606", X"25FE", X"25F5", X"25ED", X"25E4", X"25DB", 
X"25D3", X"25CA", X"25C2", X"25B9", X"25B1", X"25A8", X"25A0", X"2597", X"258F", X"2586", 
X"257E", X"2575", X"256C", X"2564", X"255B", X"2553", X"254A", X"2542", X"2539", X"2531", 
X"2528", X"251F", X"2517", X"250E", X"2506", X"24FD", X"24F5", X"24EC", X"24E4", X"24DB", 
X"24D3", X"24CA", X"24C1", X"24B9", X"24B0", X"24A8", X"249F", X"2497", X"248E", X"2485", 
X"247D", X"2474", X"246C", X"2463", X"245B", X"2452", X"2449", X"2441", X"2438", X"2430", 
X"2427", X"241F", X"2416", X"240D", X"2405", X"23FC", X"23F4", X"23EB", X"23E3", X"23DA", 
X"23D1", X"23C9", X"23C0", X"23B8", X"23AF", X"23A7", X"239E", X"2395", X"238D", X"2384", 
X"237C", X"2373", X"236A", X"2362", X"2359", X"2351", X"2348", X"233F", X"2337", X"232E", 
X"2326", X"231D", X"2315", X"230C", X"2303", X"22FB", X"22F2", X"22EA", X"22E1", X"22D8", 
X"22D0", X"22C7", X"22BF", X"22B6", X"22AD", X"22A5", X"229C", X"2294", X"228B", X"2282", 
X"227A", X"2271", X"2269", X"2260", X"2257", X"224F", X"2246", X"223D", X"2235", X"222C", 
X"2224", X"221B", X"2212", X"220A", X"2201", X"21F9", X"21F0", X"21E7", X"21DF", X"21D6", 
X"21CD", X"21C5", X"21BC", X"21B4", X"21AB", X"21A2", X"219A", X"2191", X"2189", X"2180", 
X"2177", X"216F", X"2166", X"215D", X"2155", X"214C", X"2144", X"213B", X"2132", X"212A", 
X"2121", X"2118", X"2110", X"2107", X"20FE", X"20F6", X"20ED", X"20E5", X"20DC", X"20D3", 
X"20CB", X"20C2", X"20B9", X"20B1", X"20A8", X"209F", X"2097", X"208E", X"2086", X"207D", 
X"2074", X"206C", X"2063", X"205A", X"2052", X"2049", X"2040", X"2038", X"202F", X"2026", 
X"201E", X"2015", X"200C", X"2004", X"1FFB", X"1FF2", X"1FEA", X"1FE1", X"1FD9", X"1FD0", 
X"1FC7", X"1FBF", X"1FB6", X"1FAD", X"1FA5", X"1F9C", X"1F93", X"1F8B", X"1F82", X"1F79", 
X"1F71", X"1F68", X"1F5F", X"1F57", X"1F4E", X"1F45", X"1F3D", X"1F34", X"1F2B", X"1F23", 
X"1F1A", X"1F11", X"1F09", X"1F00", X"1EF7", X"1EEF", X"1EE6", X"1EDD", X"1ED5", X"1ECC", 
X"1EC3", X"1EBB", X"1EB2", X"1EA9", X"1EA1", X"1E98", X"1E8F", X"1E87", X"1E7E", X"1E75", 
X"1E6C", X"1E64", X"1E5B", X"1E52", X"1E4A", X"1E41", X"1E38", X"1E30", X"1E27", X"1E1E", 
X"1E16", X"1E0D", X"1E04", X"1DFC", X"1DF3", X"1DEA", X"1DE2", X"1DD9", X"1DD0", X"1DC7", 
X"1DBF", X"1DB6", X"1DAD", X"1DA5", X"1D9C", X"1D93", X"1D8B", X"1D82", X"1D79", X"1D71", 
X"1D68", X"1D5F", X"1D56", X"1D4E", X"1D45", X"1D3C", X"1D34", X"1D2B", X"1D22", X"1D1A", 
X"1D11", X"1D08", X"1CFF", X"1CF7", X"1CEE", X"1CE5", X"1CDD", X"1CD4", X"1CCB", X"1CC2", 
X"1CBA", X"1CB1", X"1CA8", X"1CA0", X"1C97", X"1C8E", X"1C86", X"1C7D", X"1C74", X"1C6B", 
X"1C63", X"1C5A", X"1C51", X"1C49", X"1C40", X"1C37", X"1C2E", X"1C26", X"1C1D", X"1C14", 
X"1C0C", X"1C03", X"1BFA", X"1BF1", X"1BE9", X"1BE0", X"1BD7", X"1BCE", X"1BC6", X"1BBD", 
X"1BB4", X"1BAC", X"1BA3", X"1B9A", X"1B91", X"1B89", X"1B80", X"1B77", X"1B6E", X"1B66", 
X"1B5D", X"1B54", X"1B4C", X"1B43", X"1B3A", X"1B31", X"1B29", X"1B20", X"1B17", X"1B0E", 
X"1B06", X"1AFD", X"1AF4", X"1AEB", X"1AE3", X"1ADA", X"1AD1", X"1AC9", X"1AC0", X"1AB7", 
X"1AAE", X"1AA6", X"1A9D", X"1A94", X"1A8B", X"1A83", X"1A7A", X"1A71", X"1A68", X"1A60", 
X"1A57", X"1A4E", X"1A45", X"1A3D", X"1A34", X"1A2B", X"1A22", X"1A1A", X"1A11", X"1A08", 
X"19FF", X"19F7", X"19EE", X"19E5", X"19DC", X"19D4", X"19CB", X"19C2", X"19B9", X"19B1", 
X"19A8", X"199F", X"1996", X"198E", X"1985", X"197C", X"1973", X"196B", X"1962", X"1959", 
X"1950", X"1948", X"193F", X"1936", X"192D", X"1925", X"191C", X"1913", X"190A", X"1901", 
X"18F9", X"18F0", X"18E7", X"18DE", X"18D6", X"18CD", X"18C4", X"18BB", X"18B3", X"18AA", 
X"18A1", X"1898", X"1890", X"1887", X"187E", X"1875", X"186C", X"1864", X"185B", X"1852", 
X"1849", X"1841", X"1838", X"182F", X"1826", X"181D", X"1815", X"180C", X"1803", X"17FA", 
X"17F2", X"17E9", X"17E0", X"17D7", X"17CE", X"17C6", X"17BD", X"17B4", X"17AB", X"17A3", 
X"179A", X"1791", X"1788", X"177F", X"1777", X"176E", X"1765", X"175C", X"1753", X"174B", 
X"1742", X"1739", X"1730", X"1728", X"171F", X"1716", X"170D", X"1704", X"16FC", X"16F3", 
X"16EA", X"16E1", X"16D8", X"16D0", X"16C7", X"16BE", X"16B5", X"16AC", X"16A4", X"169B", 
X"1692", X"1689", X"1680", X"1678", X"166F", X"1666", X"165D", X"1655", X"164C", X"1643", 
X"163A", X"1631", X"1629", X"1620", X"1617", X"160E", X"1605", X"15FC", X"15F4", X"15EB", 
X"15E2", X"15D9", X"15D0", X"15C8", X"15BF", X"15B6", X"15AD", X"15A4", X"159C", X"1593", 
X"158A", X"1581", X"1578", X"1570", X"1567", X"155E", X"1555", X"154C", X"1544", X"153B", 
X"1532", X"1529", X"1520", X"1517", X"150F", X"1506", X"14FD", X"14F4", X"14EB", X"14E3", 
X"14DA", X"14D1", X"14C8", X"14BF", X"14B6", X"14AE", X"14A5", X"149C", X"1493", X"148A", 
X"1482", X"1479", X"1470", X"1467", X"145E", X"1455", X"144D", X"1444", X"143B", X"1432", 
X"1429", X"1421", X"1418", X"140F", X"1406", X"13FD", X"13F4", X"13EC", X"13E3", X"13DA", 
X"13D1", X"13C8", X"13BF", X"13B7", X"13AE", X"13A5", X"139C", X"1393", X"138A", X"1382", 
X"1379", X"1370", X"1367", X"135E", X"1355", X"134D", X"1344", X"133B", X"1332", X"1329", 
X"1320", X"1318", X"130F", X"1306", X"12FD", X"12F4", X"12EB", X"12E3", X"12DA", X"12D1", 
X"12C8", X"12BF", X"12B6", X"12AE", X"12A5", X"129C", X"1293", X"128A", X"1281", X"1278", 
X"1270", X"1267", X"125E", X"1255", X"124C", X"1243", X"123B", X"1232", X"1229", X"1220", 
X"1217", X"120E", X"1206", X"11FD", X"11F4", X"11EB", X"11E2", X"11D9", X"11D0", X"11C8", 
X"11BF", X"11B6", X"11AD", X"11A4", X"119B", X"1192", X"118A", X"1181", X"1178", X"116F", 
X"1166", X"115D", X"1155", X"114C", X"1143", X"113A", X"1131", X"1128", X"111F", X"1117", 
X"110E", X"1105", X"10FC", X"10F3", X"10EA", X"10E1", X"10D9", X"10D0", X"10C7", X"10BE", 
X"10B5", X"10AC", X"10A3", X"109B", X"1092", X"1089", X"1080", X"1077", X"106E", X"1065", 
X"105C", X"1054", X"104B", X"1042", X"1039", X"1030", X"1027", X"101E", X"1016", X"100D", 
X"1004", X"0FFB", X"0FF2", X"0FE9", X"0FE0", X"0FD7", X"0FCF", X"0FC6", X"0FBD", X"0FB4", 
X"0FAB", X"0FA2", X"0F99", X"0F91", X"0F88", X"0F7F", X"0F76", X"0F6D", X"0F64", X"0F5B", 
X"0F52", X"0F4A", X"0F41", X"0F38", X"0F2F", X"0F26", X"0F1D", X"0F14", X"0F0B", X"0F03", 
X"0EFA", X"0EF1", X"0EE8", X"0EDF", X"0ED6", X"0ECD", X"0EC4", X"0EBC", X"0EB3", X"0EAA", 
X"0EA1", X"0E98", X"0E8F", X"0E86", X"0E7D", X"0E75", X"0E6C", X"0E63", X"0E5A", X"0E51", 
X"0E48", X"0E3F", X"0E36", X"0E2E", X"0E25", X"0E1C", X"0E13", X"0E0A", X"0E01", X"0DF8", 
X"0DEF", X"0DE6", X"0DDE", X"0DD5", X"0DCC", X"0DC3", X"0DBA", X"0DB1", X"0DA8", X"0D9F", 
X"0D97", X"0D8E", X"0D85", X"0D7C", X"0D73", X"0D6A", X"0D61", X"0D58", X"0D4F", X"0D47", 
X"0D3E", X"0D35", X"0D2C", X"0D23", X"0D1A", X"0D11", X"0D08", X"0CFF", X"0CF7", X"0CEE", 
X"0CE5", X"0CDC", X"0CD3", X"0CCA", X"0CC1", X"0CB8", X"0CAF", X"0CA7", X"0C9E", X"0C95", 
X"0C8C", X"0C83", X"0C7A", X"0C71", X"0C68", X"0C5F", X"0C56", X"0C4E", X"0C45", X"0C3C", 
X"0C33", X"0C2A", X"0C21", X"0C18", X"0C0F", X"0C06", X"0BFE", X"0BF5", X"0BEC", X"0BE3", 
X"0BDA", X"0BD1", X"0BC8", X"0BBF", X"0BB6", X"0BAD", X"0BA5", X"0B9C", X"0B93", X"0B8A", 
X"0B81", X"0B78", X"0B6F", X"0B66", X"0B5D", X"0B54", X"0B4C", X"0B43", X"0B3A", X"0B31", 
X"0B28", X"0B1F", X"0B16", X"0B0D", X"0B04", X"0AFB", X"0AF3", X"0AEA", X"0AE1", X"0AD8", 
X"0ACF", X"0AC6", X"0ABD", X"0AB4", X"0AAB", X"0AA2", X"0A99", X"0A91", X"0A88", X"0A7F", 
X"0A76", X"0A6D", X"0A64", X"0A5B", X"0A52", X"0A49", X"0A40", X"0A37", X"0A2F", X"0A26", 
X"0A1D", X"0A14", X"0A0B", X"0A02", X"09F9", X"09F0", X"09E7", X"09DE", X"09D5", X"09CD", 
X"09C4", X"09BB", X"09B2", X"09A9", X"09A0", X"0997", X"098E", X"0985", X"097C", X"0973", 
X"096B", X"0962", X"0959", X"0950", X"0947", X"093E", X"0935", X"092C", X"0923", X"091A", 
X"0911", X"0909", X"0900", X"08F7", X"08EE", X"08E5", X"08DC", X"08D3", X"08CA", X"08C1", 
X"08B8", X"08AF", X"08A6", X"089E", X"0895", X"088C", X"0883", X"087A", X"0871", X"0868", 
X"085F", X"0856", X"084D", X"0844", X"083B", X"0833", X"082A", X"0821", X"0818", X"080F", 
X"0806", X"07FD", X"07F4", X"07EB", X"07E2", X"07D9", X"07D0", X"07C8", X"07BF", X"07B6", 
X"07AD", X"07A4", X"079B", X"0792", X"0789", X"0780", X"0777", X"076E", X"0765", X"075C", 
X"0754", X"074B", X"0742", X"0739", X"0730", X"0727", X"071E", X"0715", X"070C", X"0703", 
X"06FA", X"06F1", X"06E8", X"06E0", X"06D7", X"06CE", X"06C5", X"06BC", X"06B3", X"06AA", 
X"06A1", X"0698", X"068F", X"0686", X"067D", X"0674", X"066C", X"0663", X"065A", X"0651", 
X"0648", X"063F", X"0636", X"062D", X"0624", X"061B", X"0612", X"0609", X"0600", X"05F8", 
X"05EF", X"05E6", X"05DD", X"05D4", X"05CB", X"05C2", X"05B9", X"05B0", X"05A7", X"059E", 
X"0595", X"058C", X"0583", X"057B", X"0572", X"0569", X"0560", X"0557", X"054E", X"0545", 
X"053C", X"0533", X"052A", X"0521", X"0518", X"050F", X"0506", X"04FE", X"04F5", X"04EC", 
X"04E3", X"04DA", X"04D1", X"04C8", X"04BF", X"04B6", X"04AD", X"04A4", X"049B", X"0492", 
X"0489", X"0481", X"0478", X"046F", X"0466", X"045D", X"0454", X"044B", X"0442", X"0439", 
X"0430", X"0427", X"041E", X"0415", X"040C", X"0403", X"03FB", X"03F2", X"03E9", X"03E0", 
X"03D7", X"03CE", X"03C5", X"03BC", X"03B3", X"03AA", X"03A1", X"0398", X"038F", X"0386", 
X"037D", X"0375", X"036C", X"0363", X"035A", X"0351", X"0348", X"033F", X"0336", X"032D", 
X"0324", X"031B", X"0312", X"0309", X"0300", X"02F7", X"02EF", X"02E6", X"02DD", X"02D4", 
X"02CB", X"02C2", X"02B9", X"02B0", X"02A7", X"029E", X"0295", X"028C", X"0283", X"027A", 
X"0271", X"0269", X"0260", X"0257", X"024E", X"0245", X"023C", X"0233", X"022A", X"0221", 
X"0218", X"020F", X"0206", X"01FD", X"01F4", X"01EB", X"01E3", X"01DA", X"01D1", X"01C8", 
X"01BF", X"01B6", X"01AD", X"01A4", X"019B", X"0192", X"0189", X"0180", X"0177", X"016E", 
X"0165", X"015D", X"0154", X"014B", X"0142", X"0139", X"0130", X"0127", X"011E", X"0115", 
X"010C", X"0103", X"00FA", X"00F1", X"00E8", X"00DF", X"00D6", X"00CE", X"00C5", X"00BC", 
X"00B3", X"00AA", X"00A1", X"0098", X"008F", X"0086", X"007D", X"0074", X"006B", X"0062", 
X"0059", X"0050", X"0047", X"003F", X"0036", X"002D", X"0024", X"001B", X"0012", X"0009", 
X"0000", X"8009", X"8012", X"801B", X"8024", X"802D", X"8036", X"803F", X"8047", X"8050", 
X"8059", X"8062", X"806B", X"8074", X"807D", X"8086", X"808F", X"8098", X"80A1", X"80AA", 
X"80B3", X"80BC", X"80C5", X"80CE", X"80D6", X"80DF", X"80E8", X"80F1", X"80FA", X"8103", 
X"810C", X"8115", X"811E", X"8127", X"8130", X"8139", X"8142", X"814B", X"8154", X"815D", 
X"8165", X"816E", X"8177", X"8180", X"8189", X"8192", X"819B", X"81A4", X"81AD", X"81B6", 
X"81BF", X"81C8", X"81D1", X"81DA", X"81E3", X"81EB", X"81F4", X"81FD", X"8206", X"820F", 
X"8218", X"8221", X"822A", X"8233", X"823C", X"8245", X"824E", X"8257", X"8260", X"8269", 
X"8271", X"827A", X"8283", X"828C", X"8295", X"829E", X"82A7", X"82B0", X"82B9", X"82C2", 
X"82CB", X"82D4", X"82DD", X"82E6", X"82EF", X"82F7", X"8300", X"8309", X"8312", X"831B", 
X"8324", X"832D", X"8336", X"833F", X"8348", X"8351", X"835A", X"8363", X"836C", X"8375", 
X"837D", X"8386", X"838F", X"8398", X"83A1", X"83AA", X"83B3", X"83BC", X"83C5", X"83CE", 
X"83D7", X"83E0", X"83E9", X"83F2", X"83FB", X"8403", X"840C", X"8415", X"841E", X"8427", 
X"8430", X"8439", X"8442", X"844B", X"8454", X"845D", X"8466", X"846F", X"8478", X"8481", 
X"8489", X"8492", X"849B", X"84A4", X"84AD", X"84B6", X"84BF", X"84C8", X"84D1", X"84DA", 
X"84E3", X"84EC", X"84F5", X"84FE", X"8506", X"850F", X"8518", X"8521", X"852A", X"8533", 
X"853C", X"8545", X"854E", X"8557", X"8560", X"8569", X"8572", X"857B", X"8583", X"858C", 
X"8595", X"859E", X"85A7", X"85B0", X"85B9", X"85C2", X"85CB", X"85D4", X"85DD", X"85E6", 
X"85EF", X"85F8", X"8600", X"8609", X"8612", X"861B", X"8624", X"862D", X"8636", X"863F", 
X"8648", X"8651", X"865A", X"8663", X"866C", X"8674", X"867D", X"8686", X"868F", X"8698", 
X"86A1", X"86AA", X"86B3", X"86BC", X"86C5", X"86CE", X"86D7", X"86E0", X"86E8", X"86F1", 
X"86FA", X"8703", X"870C", X"8715", X"871E", X"8727", X"8730", X"8739", X"8742", X"874B", 
X"8754", X"875C", X"8765", X"876E", X"8777", X"8780", X"8789", X"8792", X"879B", X"87A4", 
X"87AD", X"87B6", X"87BF", X"87C8", X"87D0", X"87D9", X"87E2", X"87EB", X"87F4", X"87FD", 
X"8806", X"880F", X"8818", X"8821", X"882A", X"8833", X"883B", X"8844", X"884D", X"8856", 
X"885F", X"8868", X"8871", X"887A", X"8883", X"888C", X"8895", X"889E", X"88A6", X"88AF", 
X"88B8", X"88C1", X"88CA", X"88D3", X"88DC", X"88E5", X"88EE", X"88F7", X"8900", X"8909", 
X"8911", X"891A", X"8923", X"892C", X"8935", X"893E", X"8947", X"8950", X"8959", X"8962", 
X"896B", X"8973", X"897C", X"8985", X"898E", X"8997", X"89A0", X"89A9", X"89B2", X"89BB", 
X"89C4", X"89CD", X"89D5", X"89DE", X"89E7", X"89F0", X"89F9", X"8A02", X"8A0B", X"8A14", 
X"8A1D", X"8A26", X"8A2F", X"8A37", X"8A40", X"8A49", X"8A52", X"8A5B", X"8A64", X"8A6D", 
X"8A76", X"8A7F", X"8A88", X"8A91", X"8A99", X"8AA2", X"8AAB", X"8AB4", X"8ABD", X"8AC6", 
X"8ACF", X"8AD8", X"8AE1", X"8AEA", X"8AF3", X"8AFB", X"8B04", X"8B0D", X"8B16", X"8B1F", 
X"8B28", X"8B31", X"8B3A", X"8B43", X"8B4C", X"8B54", X"8B5D", X"8B66", X"8B6F", X"8B78", 
X"8B81", X"8B8A", X"8B93", X"8B9C", X"8BA5", X"8BAD", X"8BB6", X"8BBF", X"8BC8", X"8BD1", 
X"8BDA", X"8BE3", X"8BEC", X"8BF5", X"8BFE", X"8C06", X"8C0F", X"8C18", X"8C21", X"8C2A", 
X"8C33", X"8C3C", X"8C45", X"8C4E", X"8C56", X"8C5F", X"8C68", X"8C71", X"8C7A", X"8C83", 
X"8C8C", X"8C95", X"8C9E", X"8CA7", X"8CAF", X"8CB8", X"8CC1", X"8CCA", X"8CD3", X"8CDC", 
X"8CE5", X"8CEE", X"8CF7", X"8CFF", X"8D08", X"8D11", X"8D1A", X"8D23", X"8D2C", X"8D35", 
X"8D3E", X"8D47", X"8D4F", X"8D58", X"8D61", X"8D6A", X"8D73", X"8D7C", X"8D85", X"8D8E", 
X"8D97", X"8D9F", X"8DA8", X"8DB1", X"8DBA", X"8DC3", X"8DCC", X"8DD5", X"8DDE", X"8DE6", 
X"8DEF", X"8DF8", X"8E01", X"8E0A", X"8E13", X"8E1C", X"8E25", X"8E2E", X"8E36", X"8E3F", 
X"8E48", X"8E51", X"8E5A", X"8E63", X"8E6C", X"8E75", X"8E7D", X"8E86", X"8E8F", X"8E98", 
X"8EA1", X"8EAA", X"8EB3", X"8EBC", X"8EC4", X"8ECD", X"8ED6", X"8EDF", X"8EE8", X"8EF1", 
X"8EFA", X"8F03", X"8F0B", X"8F14", X"8F1D", X"8F26", X"8F2F", X"8F38", X"8F41", X"8F4A", 
X"8F52", X"8F5B", X"8F64", X"8F6D", X"8F76", X"8F7F", X"8F88", X"8F91", X"8F99", X"8FA2", 
X"8FAB", X"8FB4", X"8FBD", X"8FC6", X"8FCF", X"8FD7", X"8FE0", X"8FE9", X"8FF2", X"8FFB", 
X"9004", X"900D", X"9016", X"901E", X"9027", X"9030", X"9039", X"9042", X"904B", X"9054", 
X"905C", X"9065", X"906E", X"9077", X"9080", X"9089", X"9092", X"909B", X"90A3", X"90AC", 
X"90B5", X"90BE", X"90C7", X"90D0", X"90D9", X"90E1", X"90EA", X"90F3", X"90FC", X"9105", 
X"910E", X"9117", X"911F", X"9128", X"9131", X"913A", X"9143", X"914C", X"9155", X"915D", 
X"9166", X"916F", X"9178", X"9181", X"918A", X"9192", X"919B", X"91A4", X"91AD", X"91B6", 
X"91BF", X"91C8", X"91D0", X"91D9", X"91E2", X"91EB", X"91F4", X"91FD", X"9206", X"920E", 
X"9217", X"9220", X"9229", X"9232", X"923B", X"9243", X"924C", X"9255", X"925E", X"9267", 
X"9270", X"9278", X"9281", X"928A", X"9293", X"929C", X"92A5", X"92AE", X"92B6", X"92BF", 
X"92C8", X"92D1", X"92DA", X"92E3", X"92EB", X"92F4", X"92FD", X"9306", X"930F", X"9318", 
X"9320", X"9329", X"9332", X"933B", X"9344", X"934D", X"9355", X"935E", X"9367", X"9370", 
X"9379", X"9382", X"938A", X"9393", X"939C", X"93A5", X"93AE", X"93B7", X"93BF", X"93C8", 
X"93D1", X"93DA", X"93E3", X"93EC", X"93F4", X"93FD", X"9406", X"940F", X"9418", X"9421", 
X"9429", X"9432", X"943B", X"9444", X"944D", X"9455", X"945E", X"9467", X"9470", X"9479", 
X"9482", X"948A", X"9493", X"949C", X"94A5", X"94AE", X"94B6", X"94BF", X"94C8", X"94D1", 
X"94DA", X"94E3", X"94EB", X"94F4", X"94FD", X"9506", X"950F", X"9517", X"9520", X"9529", 
X"9532", X"953B", X"9544", X"954C", X"9555", X"955E", X"9567", X"9570", X"9578", X"9581", 
X"958A", X"9593", X"959C", X"95A4", X"95AD", X"95B6", X"95BF", X"95C8", X"95D0", X"95D9", 
X"95E2", X"95EB", X"95F4", X"95FC", X"9605", X"960E", X"9617", X"9620", X"9629", X"9631", 
X"963A", X"9643", X"964C", X"9655", X"965D", X"9666", X"966F", X"9678", X"9680", X"9689", 
X"9692", X"969B", X"96A4", X"96AC", X"96B5", X"96BE", X"96C7", X"96D0", X"96D8", X"96E1", 
X"96EA", X"96F3", X"96FC", X"9704", X"970D", X"9716", X"971F", X"9728", X"9730", X"9739", 
X"9742", X"974B", X"9753", X"975C", X"9765", X"976E", X"9777", X"977F", X"9788", X"9791", 
X"979A", X"97A3", X"97AB", X"97B4", X"97BD", X"97C6", X"97CE", X"97D7", X"97E0", X"97E9", 
X"97F2", X"97FA", X"9803", X"980C", X"9815", X"981D", X"9826", X"982F", X"9838", X"9841", 
X"9849", X"9852", X"985B", X"9864", X"986C", X"9875", X"987E", X"9887", X"9890", X"9898", 
X"98A1", X"98AA", X"98B3", X"98BB", X"98C4", X"98CD", X"98D6", X"98DE", X"98E7", X"98F0", 
X"98F9", X"9901", X"990A", X"9913", X"991C", X"9925", X"992D", X"9936", X"993F", X"9948", 
X"9950", X"9959", X"9962", X"996B", X"9973", X"997C", X"9985", X"998E", X"9996", X"999F", 
X"99A8", X"99B1", X"99B9", X"99C2", X"99CB", X"99D4", X"99DC", X"99E5", X"99EE", X"99F7", 
X"99FF", X"9A08", X"9A11", X"9A1A", X"9A22", X"9A2B", X"9A34", X"9A3D", X"9A45", X"9A4E", 
X"9A57", X"9A60", X"9A68", X"9A71", X"9A7A", X"9A83", X"9A8B", X"9A94", X"9A9D", X"9AA6", 
X"9AAE", X"9AB7", X"9AC0", X"9AC9", X"9AD1", X"9ADA", X"9AE3", X"9AEB", X"9AF4", X"9AFD", 
X"9B06", X"9B0E", X"9B17", X"9B20", X"9B29", X"9B31", X"9B3A", X"9B43", X"9B4C", X"9B54", 
X"9B5D", X"9B66", X"9B6E", X"9B77", X"9B80", X"9B89", X"9B91", X"9B9A", X"9BA3", X"9BAC", 
X"9BB4", X"9BBD", X"9BC6", X"9BCE", X"9BD7", X"9BE0", X"9BE9", X"9BF1", X"9BFA", X"9C03", 
X"9C0C", X"9C14", X"9C1D", X"9C26", X"9C2E", X"9C37", X"9C40", X"9C49", X"9C51", X"9C5A", 
X"9C63", X"9C6B", X"9C74", X"9C7D", X"9C86", X"9C8E", X"9C97", X"9CA0", X"9CA8", X"9CB1", 
X"9CBA", X"9CC2", X"9CCB", X"9CD4", X"9CDD", X"9CE5", X"9CEE", X"9CF7", X"9CFF", X"9D08", 
X"9D11", X"9D1A", X"9D22", X"9D2B", X"9D34", X"9D3C", X"9D45", X"9D4E", X"9D56", X"9D5F", 
X"9D68", X"9D71", X"9D79", X"9D82", X"9D8B", X"9D93", X"9D9C", X"9DA5", X"9DAD", X"9DB6", 
X"9DBF", X"9DC7", X"9DD0", X"9DD9", X"9DE2", X"9DEA", X"9DF3", X"9DFC", X"9E04", X"9E0D", 
X"9E16", X"9E1E", X"9E27", X"9E30", X"9E38", X"9E41", X"9E4A", X"9E52", X"9E5B", X"9E64", 
X"9E6C", X"9E75", X"9E7E", X"9E87", X"9E8F", X"9E98", X"9EA1", X"9EA9", X"9EB2", X"9EBB", 
X"9EC3", X"9ECC", X"9ED5", X"9EDD", X"9EE6", X"9EEF", X"9EF7", X"9F00", X"9F09", X"9F11", 
X"9F1A", X"9F23", X"9F2B", X"9F34", X"9F3D", X"9F45", X"9F4E", X"9F57", X"9F5F", X"9F68", 
X"9F71", X"9F79", X"9F82", X"9F8B", X"9F93", X"9F9C", X"9FA5", X"9FAD", X"9FB6", X"9FBF", 
X"9FC7", X"9FD0", X"9FD9", X"9FE1", X"9FEA", X"9FF2", X"9FFB", X"A004", X"A00C", X"A015", 
X"A01E", X"A026", X"A02F", X"A038", X"A040", X"A049", X"A052", X"A05A", X"A063", X"A06C", 
X"A074", X"A07D", X"A086", X"A08E", X"A097", X"A09F", X"A0A8", X"A0B1", X"A0B9", X"A0C2", 
X"A0CB", X"A0D3", X"A0DC", X"A0E5", X"A0ED", X"A0F6", X"A0FE", X"A107", X"A110", X"A118", 
X"A121", X"A12A", X"A132", X"A13B", X"A144", X"A14C", X"A155", X"A15D", X"A166", X"A16F", 
X"A177", X"A180", X"A189", X"A191", X"A19A", X"A1A2", X"A1AB", X"A1B4", X"A1BC", X"A1C5", 
X"A1CD", X"A1D6", X"A1DF", X"A1E7", X"A1F0", X"A1F9", X"A201", X"A20A", X"A212", X"A21B", 
X"A224", X"A22C", X"A235", X"A23D", X"A246", X"A24F", X"A257", X"A260", X"A269", X"A271", 
X"A27A", X"A282", X"A28B", X"A294", X"A29C", X"A2A5", X"A2AD", X"A2B6", X"A2BF", X"A2C7", 
X"A2D0", X"A2D8", X"A2E1", X"A2EA", X"A2F2", X"A2FB", X"A303", X"A30C", X"A315", X"A31D", 
X"A326", X"A32E", X"A337", X"A33F", X"A348", X"A351", X"A359", X"A362", X"A36A", X"A373", 
X"A37C", X"A384", X"A38D", X"A395", X"A39E", X"A3A7", X"A3AF", X"A3B8", X"A3C0", X"A3C9", 
X"A3D1", X"A3DA", X"A3E3", X"A3EB", X"A3F4", X"A3FC", X"A405", X"A40D", X"A416", X"A41F", 
X"A427", X"A430", X"A438", X"A441", X"A449", X"A452", X"A45B", X"A463", X"A46C", X"A474", 
X"A47D", X"A485", X"A48E", X"A497", X"A49F", X"A4A8", X"A4B0", X"A4B9", X"A4C1", X"A4CA", 
X"A4D3", X"A4DB", X"A4E4", X"A4EC", X"A4F5", X"A4FD", X"A506", X"A50E", X"A517", X"A51F", 
X"A528", X"A531", X"A539", X"A542", X"A54A", X"A553", X"A55B", X"A564", X"A56C", X"A575", 
X"A57E", X"A586", X"A58F", X"A597", X"A5A0", X"A5A8", X"A5B1", X"A5B9", X"A5C2", X"A5CA", 
X"A5D3", X"A5DB", X"A5E4", X"A5ED", X"A5F5", X"A5FE", X"A606", X"A60F", X"A617", X"A620", 
X"A628", X"A631", X"A639", X"A642", X"A64A", X"A653", X"A65B", X"A664", X"A66C", X"A675", 
X"A67E", X"A686", X"A68F", X"A697", X"A6A0", X"A6A8", X"A6B1", X"A6B9", X"A6C2", X"A6CA", 
X"A6D3", X"A6DB", X"A6E4", X"A6EC", X"A6F5", X"A6FD", X"A706", X"A70E", X"A717", X"A71F", 
X"A728", X"A730", X"A739", X"A741", X"A74A", X"A752", X"A75B", X"A763", X"A76C", X"A774", 
X"A77D", X"A785", X"A78E", X"A796", X"A79F", X"A7A7", X"A7B0", X"A7B8", X"A7C1", X"A7C9", 
X"A7D2", X"A7DA", X"A7E3", X"A7EB", X"A7F4", X"A7FC", X"A805", X"A80D", X"A816", X"A81E", 
X"A827", X"A82F", X"A838", X"A840", X"A849", X"A851", X"A85A", X"A862", X"A86B", X"A873", 
X"A87C", X"A884", X"A88C", X"A895", X"A89D", X"A8A6", X"A8AE", X"A8B7", X"A8BF", X"A8C8", 
X"A8D0", X"A8D9", X"A8E1", X"A8EA", X"A8F2", X"A8FB", X"A903", X"A90C", X"A914", X"A91C", 
X"A925", X"A92D", X"A936", X"A93E", X"A947", X"A94F", X"A958", X"A960", X"A969", X"A971", 
X"A97A", X"A982", X"A98A", X"A993", X"A99B", X"A9A4", X"A9AC", X"A9B5", X"A9BD", X"A9C6", 
X"A9CE", X"A9D6", X"A9DF", X"A9E7", X"A9F0", X"A9F8", X"AA01", X"AA09", X"AA12", X"AA1A", 
X"AA22", X"AA2B", X"AA33", X"AA3C", X"AA44", X"AA4D", X"AA55", X"AA5D", X"AA66", X"AA6E", 
X"AA77", X"AA7F", X"AA88", X"AA90", X"AA98", X"AAA1", X"AAA9", X"AAB2", X"AABA", X"AAC3", 
X"AACB", X"AAD3", X"AADC", X"AAE4", X"AAED", X"AAF5", X"AAFE", X"AB06", X"AB0E", X"AB17", 
X"AB1F", X"AB28", X"AB30", X"AB38", X"AB41", X"AB49", X"AB52", X"AB5A", X"AB62", X"AB6B", 
X"AB73", X"AB7C", X"AB84", X"AB8D", X"AB95", X"AB9D", X"ABA6", X"ABAE", X"ABB7", X"ABBF", 
X"ABC7", X"ABD0", X"ABD8", X"ABE1", X"ABE9", X"ABF1", X"ABFA", X"AC02", X"AC0A", X"AC13", 
X"AC1B", X"AC24", X"AC2C", X"AC34", X"AC3D", X"AC45", X"AC4E", X"AC56", X"AC5E", X"AC67", 
X"AC6F", X"AC77", X"AC80", X"AC88", X"AC91", X"AC99", X"ACA1", X"ACAA", X"ACB2", X"ACBA", 
X"ACC3", X"ACCB", X"ACD4", X"ACDC", X"ACE4", X"ACED", X"ACF5", X"ACFD", X"AD06", X"AD0E", 
X"AD17", X"AD1F", X"AD27", X"AD30", X"AD38", X"AD40", X"AD49", X"AD51", X"AD59", X"AD62", 
X"AD6A", X"AD72", X"AD7B", X"AD83", X"AD8C", X"AD94", X"AD9C", X"ADA5", X"ADAD", X"ADB5", 
X"ADBE", X"ADC6", X"ADCE", X"ADD7", X"ADDF", X"ADE7", X"ADF0", X"ADF8", X"AE00", X"AE09", 
X"AE11", X"AE19", X"AE22", X"AE2A", X"AE32", X"AE3B", X"AE43", X"AE4B", X"AE54", X"AE5C", 
X"AE64", X"AE6D", X"AE75", X"AE7D", X"AE86", X"AE8E", X"AE96", X"AE9F", X"AEA7", X"AEAF", 
X"AEB8", X"AEC0", X"AEC8", X"AED1", X"AED9", X"AEE1", X"AEEA", X"AEF2", X"AEFA", X"AF02", 
X"AF0B", X"AF13", X"AF1B", X"AF24", X"AF2C", X"AF34", X"AF3D", X"AF45", X"AF4D", X"AF56", 
X"AF5E", X"AF66", X"AF6E", X"AF77", X"AF7F", X"AF87", X"AF90", X"AF98", X"AFA0", X"AFA9", 
X"AFB1", X"AFB9", X"AFC1", X"AFCA", X"AFD2", X"AFDA", X"AFE3", X"AFEB", X"AFF3", X"AFFB", 
X"B004", X"B00C", X"B014", X"B01D", X"B025", X"B02D", X"B035", X"B03E", X"B046", X"B04E", 
X"B056", X"B05F", X"B067", X"B06F", X"B078", X"B080", X"B088", X"B090", X"B099", X"B0A1", 
X"B0A9", X"B0B1", X"B0BA", X"B0C2", X"B0CA", X"B0D2", X"B0DB", X"B0E3", X"B0EB", X"B0F4", 
X"B0FC", X"B104", X"B10C", X"B115", X"B11D", X"B125", X"B12D", X"B136", X"B13E", X"B146", 
X"B14E", X"B157", X"B15F", X"B167", X"B16F", X"B178", X"B180", X"B188", X"B190", X"B198", 
X"B1A1", X"B1A9", X"B1B1", X"B1B9", X"B1C2", X"B1CA", X"B1D2", X"B1DA", X"B1E3", X"B1EB", 
X"B1F3", X"B1FB", X"B203", X"B20C", X"B214", X"B21C", X"B224", X"B22D", X"B235", X"B23D", 
X"B245", X"B24D", X"B256", X"B25E", X"B266", X"B26E", X"B277", X"B27F", X"B287", X"B28F", 
X"B297", X"B2A0", X"B2A8", X"B2B0", X"B2B8", X"B2C0", X"B2C9", X"B2D1", X"B2D9", X"B2E1", 
X"B2E9", X"B2F2", X"B2FA", X"B302", X"B30A", X"B312", X"B31B", X"B323", X"B32B", X"B333", 
X"B33B", X"B344", X"B34C", X"B354", X"B35C", X"B364", X"B36C", X"B375", X"B37D", X"B385", 
X"B38D", X"B395", X"B39E", X"B3A6", X"B3AE", X"B3B6", X"B3BE", X"B3C6", X"B3CF", X"B3D7", 
X"B3DF", X"B3E7", X"B3EF", X"B3F7", X"B400", X"B408", X"B410", X"B418", X"B420", X"B428", 
X"B431", X"B439", X"B441", X"B449", X"B451", X"B459", X"B462", X"B46A", X"B472", X"B47A", 
X"B482", X"B48A", X"B492", X"B49B", X"B4A3", X"B4AB", X"B4B3", X"B4BB", X"B4C3", X"B4CB", 
X"B4D4", X"B4DC", X"B4E4", X"B4EC", X"B4F4", X"B4FC", X"B504", X"B50D", X"B515", X"B51D", 
X"B525", X"B52D", X"B535", X"B53D", X"B545", X"B54E", X"B556", X"B55E", X"B566", X"B56E", 
X"B576", X"B57E", X"B586", X"B58F", X"B597", X"B59F", X"B5A7", X"B5AF", X"B5B7", X"B5BF", 
X"B5C7", X"B5CF", X"B5D8", X"B5E0", X"B5E8", X"B5F0", X"B5F8", X"B600", X"B608", X"B610", 
X"B618", X"B620", X"B629", X"B631", X"B639", X"B641", X"B649", X"B651", X"B659", X"B661", 
X"B669", X"B671", X"B679", X"B682", X"B68A", X"B692", X"B69A", X"B6A2", X"B6AA", X"B6B2", 
X"B6BA", X"B6C2", X"B6CA", X"B6D2", X"B6DA", X"B6E3", X"B6EB", X"B6F3", X"B6FB", X"B703", 
X"B70B", X"B713", X"B71B", X"B723", X"B72B", X"B733", X"B73B", X"B743", X"B74B", X"B753", 
X"B75B", X"B764", X"B76C", X"B774", X"B77C", X"B784", X"B78C", X"B794", X"B79C", X"B7A4", 
X"B7AC", X"B7B4", X"B7BC", X"B7C4", X"B7CC", X"B7D4", X"B7DC", X"B7E4", X"B7EC", X"B7F4", 
X"B7FC", X"B804", X"B80C", X"B815", X"B81D", X"B825", X"B82D", X"B835", X"B83D", X"B845", 
X"B84D", X"B855", X"B85D", X"B865", X"B86D", X"B875", X"B87D", X"B885", X"B88D", X"B895", 
X"B89D", X"B8A5", X"B8AD", X"B8B5", X"B8BD", X"B8C5", X"B8CD", X"B8D5", X"B8DD", X"B8E5", 
X"B8ED", X"B8F5", X"B8FD", X"B905", X"B90D", X"B915", X"B91D", X"B925", X"B92D", X"B935", 
X"B93D", X"B945", X"B94D", X"B955", X"B95D", X"B965", X"B96D", X"B975", X"B97D", X"B985", 
X"B98D", X"B995", X"B99D", X"B9A5", X"B9AD", X"B9B5", X"B9BD", X"B9C5", X"B9CD", X"B9D5", 
X"B9DD", X"B9E5", X"B9ED", X"B9F5", X"B9FD", X"BA04", X"BA0C", X"BA14", X"BA1C", X"BA24", 
X"BA2C", X"BA34", X"BA3C", X"BA44", X"BA4C", X"BA54", X"BA5C", X"BA64", X"BA6C", X"BA74", 
X"BA7C", X"BA84", X"BA8C", X"BA94", X"BA9C", X"BAA4", X"BAAB", X"BAB3", X"BABB", X"BAC3", 
X"BACB", X"BAD3", X"BADB", X"BAE3", X"BAEB", X"BAF3", X"BAFB", X"BB03", X"BB0B", X"BB13", 
X"BB1B", X"BB23", X"BB2A", X"BB32", X"BB3A", X"BB42", X"BB4A", X"BB52", X"BB5A", X"BB62", 
X"BB6A", X"BB72", X"BB7A", X"BB82", X"BB89", X"BB91", X"BB99", X"BBA1", X"BBA9", X"BBB1", 
X"BBB9", X"BBC1", X"BBC9", X"BBD1", X"BBD8", X"BBE0", X"BBE8", X"BBF0", X"BBF8", X"BC00", 
X"BC08", X"BC10", X"BC18", X"BC20", X"BC27", X"BC2F", X"BC37", X"BC3F", X"BC47", X"BC4F", 
X"BC57", X"BC5F", X"BC66", X"BC6E", X"BC76", X"BC7E", X"BC86", X"BC8E", X"BC96", X"BC9E", 
X"BCA5", X"BCAD", X"BCB5", X"BCBD", X"BCC5", X"BCCD", X"BCD5", X"BCDD", X"BCE4", X"BCEC", 
X"BCF4", X"BCFC", X"BD04", X"BD0C", X"BD14", X"BD1B", X"BD23", X"BD2B", X"BD33", X"BD3B", 
X"BD43", X"BD4A", X"BD52", X"BD5A", X"BD62", X"BD6A", X"BD72", X"BD7A", X"BD81", X"BD89", 
X"BD91", X"BD99", X"BDA1", X"BDA9", X"BDB0", X"BDB8", X"BDC0", X"BDC8", X"BDD0", X"BDD8", 
X"BDDF", X"BDE7", X"BDEF", X"BDF7", X"BDFF", X"BE06", X"BE0E", X"BE16", X"BE1E", X"BE26", 
X"BE2D", X"BE35", X"BE3D", X"BE45", X"BE4D", X"BE55", X"BE5C", X"BE64", X"BE6C", X"BE74", 
X"BE7C", X"BE83", X"BE8B", X"BE93", X"BE9B", X"BEA3", X"BEAA", X"BEB2", X"BEBA", X"BEC2", 
X"BEC9", X"BED1", X"BED9", X"BEE1", X"BEE9", X"BEF0", X"BEF8", X"BF00", X"BF08", X"BF10", 
X"BF17", X"BF1F", X"BF27", X"BF2F", X"BF36", X"BF3E", X"BF46", X"BF4E", X"BF55", X"BF5D", 
X"BF65", X"BF6D", X"BF75", X"BF7C", X"BF84", X"BF8C", X"BF94", X"BF9B", X"BFA3", X"BFAB", 
X"BFB3", X"BFBA", X"BFC2", X"BFCA", X"BFD2", X"BFD9", X"BFE1", X"BFE9", X"BFF1", X"BFF8", 
X"C000", X"C008", X"C00F", X"C017", X"C01F", X"C027", X"C02E", X"C036", X"C03E", X"C046", 
X"C04D", X"C055", X"C05D", X"C065", X"C06C", X"C074", X"C07C", X"C083", X"C08B", X"C093", 
X"C09B", X"C0A2", X"C0AA", X"C0B2", X"C0B9", X"C0C1", X"C0C9", X"C0D1", X"C0D8", X"C0E0", 
X"C0E8", X"C0EF", X"C0F7", X"C0FF", X"C106", X"C10E", X"C116", X"C11E", X"C125", X"C12D", 
X"C135", X"C13C", X"C144", X"C14C", X"C153", X"C15B", X"C163", X"C16A", X"C172", X"C17A", 
X"C181", X"C189", X"C191", X"C198", X"C1A0", X"C1A8", X"C1AF", X"C1B7", X"C1BF", X"C1C6", 
X"C1CE", X"C1D6", X"C1DD", X"C1E5", X"C1ED", X"C1F4", X"C1FC", X"C204", X"C20B", X"C213", 
X"C21B", X"C222", X"C22A", X"C232", X"C239", X"C241", X"C249", X"C250", X"C258", X"C260", 
X"C267", X"C26F", X"C276", X"C27E", X"C286", X"C28D", X"C295", X"C29D", X"C2A4", X"C2AC", 
X"C2B3", X"C2BB", X"C2C3", X"C2CA", X"C2D2", X"C2DA", X"C2E1", X"C2E9", X"C2F0", X"C2F8", 
X"C300", X"C307", X"C30F", X"C317", X"C31E", X"C326", X"C32D", X"C335", X"C33D", X"C344", 
X"C34C", X"C353", X"C35B", X"C363", X"C36A", X"C372", X"C379", X"C381", X"C389", X"C390", 
X"C398", X"C39F", X"C3A7", X"C3AE", X"C3B6", X"C3BE", X"C3C5", X"C3CD", X"C3D4", X"C3DC", 
X"C3E4", X"C3EB", X"C3F3", X"C3FA", X"C402", X"C409", X"C411", X"C419", X"C420", X"C428", 
X"C42F", X"C437", X"C43E", X"C446", X"C44D", X"C455", X"C45D", X"C464", X"C46C", X"C473", 
X"C47B", X"C482", X"C48A", X"C491", X"C499", X"C4A1", X"C4A8", X"C4B0", X"C4B7", X"C4BF", 
X"C4C6", X"C4CE", X"C4D5", X"C4DD", X"C4E4", X"C4EC", X"C4F3", X"C4FB", X"C502", X"C50A", 
X"C512", X"C519", X"C521", X"C528", X"C530", X"C537", X"C53F", X"C546", X"C54E", X"C555", 
X"C55D", X"C564", X"C56C", X"C573", X"C57B", X"C582", X"C58A", X"C591", X"C599", X"C5A0", 
X"C5A8", X"C5AF", X"C5B7", X"C5BE", X"C5C6", X"C5CD", X"C5D5", X"C5DC", X"C5E4", X"C5EB", 
X"C5F3", X"C5FA", X"C602", X"C609", X"C611", X"C618", X"C620", X"C627", X"C62E", X"C636", 
X"C63D", X"C645", X"C64C", X"C654", X"C65B", X"C663", X"C66A", X"C672", X"C679", X"C681", 
X"C688", X"C690", X"C697", X"C69E", X"C6A6", X"C6AD", X"C6B5", X"C6BC", X"C6C4", X"C6CB", 
X"C6D3", X"C6DA", X"C6E1", X"C6E9", X"C6F0", X"C6F8", X"C6FF", X"C707", X"C70E", X"C715", 
X"C71D", X"C724", X"C72C", X"C733", X"C73B", X"C742", X"C749", X"C751", X"C758", X"C760", 
X"C767", X"C76F", X"C776", X"C77D", X"C785", X"C78C", X"C794", X"C79B", X"C7A2", X"C7AA", 
X"C7B1", X"C7B9", X"C7C0", X"C7C7", X"C7CF", X"C7D6", X"C7DE", X"C7E5", X"C7EC", X"C7F4", 
X"C7FB", X"C803", X"C80A", X"C811", X"C819", X"C820", X"C828", X"C82F", X"C836", X"C83E", 
X"C845", X"C84C", X"C854", X"C85B", X"C863", X"C86A", X"C871", X"C879", X"C880", X"C887", 
X"C88F", X"C896", X"C89D", X"C8A5", X"C8AC", X"C8B4", X"C8BB", X"C8C2", X"C8CA", X"C8D1", 
X"C8D8", X"C8E0", X"C8E7", X"C8EE", X"C8F6", X"C8FD", X"C904", X"C90C", X"C913", X"C91A", 
X"C922", X"C929", X"C930", X"C938", X"C93F", X"C946", X"C94E", X"C955", X"C95C", X"C964", 
X"C96B", X"C972", X"C97A", X"C981", X"C988", X"C990", X"C997", X"C99E", X"C9A5", X"C9AD", 
X"C9B4", X"C9BB", X"C9C3", X"C9CA", X"C9D1", X"C9D9", X"C9E0", X"C9E7", X"C9EE", X"C9F6", 
X"C9FD", X"CA04", X"CA0C", X"CA13", X"CA1A", X"CA22", X"CA29", X"CA30", X"CA37", X"CA3F", 
X"CA46", X"CA4D", X"CA54", X"CA5C", X"CA63", X"CA6A", X"CA72", X"CA79", X"CA80", X"CA87", 
X"CA8F", X"CA96", X"CA9D", X"CAA4", X"CAAC", X"CAB3", X"CABA", X"CAC1", X"CAC9", X"CAD0", 
X"CAD7", X"CADE", X"CAE6", X"CAED", X"CAF4", X"CAFB", X"CB03", X"CB0A", X"CB11", X"CB18", 
X"CB20", X"CB27", X"CB2E", X"CB35", X"CB3D", X"CB44", X"CB4B", X"CB52", X"CB59", X"CB61", 
X"CB68", X"CB6F", X"CB76", X"CB7E", X"CB85", X"CB8C", X"CB93", X"CB9A", X"CBA2", X"CBA9", 
X"CBB0", X"CBB7", X"CBBE", X"CBC6", X"CBCD", X"CBD4", X"CBDB", X"CBE2", X"CBEA", X"CBF1", 
X"CBF8", X"CBFF", X"CC06", X"CC0E", X"CC15", X"CC1C", X"CC23", X"CC2A", X"CC32", X"CC39", 
X"CC40", X"CC47", X"CC4E", X"CC55", X"CC5D", X"CC64", X"CC6B", X"CC72", X"CC79", X"CC80", 
X"CC88", X"CC8F", X"CC96", X"CC9D", X"CCA4", X"CCAB", X"CCB3", X"CCBA", X"CCC1", X"CCC8", 
X"CCCF", X"CCD6", X"CCDD", X"CCE5", X"CCEC", X"CCF3", X"CCFA", X"CD01", X"CD08", X"CD0F", 
X"CD17", X"CD1E", X"CD25", X"CD2C", X"CD33", X"CD3A", X"CD41", X"CD48", X"CD50", X"CD57", 
X"CD5E", X"CD65", X"CD6C", X"CD73", X"CD7A", X"CD81", X"CD88", X"CD90", X"CD97", X"CD9E", 
X"CDA5", X"CDAC", X"CDB3", X"CDBA", X"CDC1", X"CDC8", X"CDD0", X"CDD7", X"CDDE", X"CDE5", 
X"CDEC", X"CDF3", X"CDFA", X"CE01", X"CE08", X"CE0F", X"CE16", X"CE1D", X"CE25", X"CE2C", 
X"CE33", X"CE3A", X"CE41", X"CE48", X"CE4F", X"CE56", X"CE5D", X"CE64", X"CE6B", X"CE72", 
X"CE79", X"CE80", X"CE88", X"CE8F", X"CE96", X"CE9D", X"CEA4", X"CEAB", X"CEB2", X"CEB9", 
X"CEC0", X"CEC7", X"CECE", X"CED5", X"CEDC", X"CEE3", X"CEEA", X"CEF1", X"CEF8", X"CEFF", 
X"CF06", X"CF0D", X"CF14", X"CF1B", X"CF22", X"CF29", X"CF30", X"CF37", X"CF3E", X"CF45", 
X"CF4D", X"CF54", X"CF5B", X"CF62", X"CF69", X"CF70", X"CF77", X"CF7E", X"CF85", X"CF8C", 
X"CF93", X"CF9A", X"CFA1", X"CFA8", X"CFAF", X"CFB6", X"CFBD", X"CFC4", X"CFCB", X"CFD2", 
X"CFD8", X"CFDF", X"CFE6", X"CFED", X"CFF4", X"CFFB", X"D002", X"D009", X"D010", X"D017", 
X"D01E", X"D025", X"D02C", X"D033", X"D03A", X"D041", X"D048", X"D04F", X"D056", X"D05D", 
X"D064", X"D06B", X"D072", X"D079", X"D080", X"D087", X"D08E", X"D095", X"D09B", X"D0A2", 
X"D0A9", X"D0B0", X"D0B7", X"D0BE", X"D0C5", X"D0CC", X"D0D3", X"D0DA", X"D0E1", X"D0E8", 
X"D0EF", X"D0F6", X"D0FC", X"D103", X"D10A", X"D111", X"D118", X"D11F", X"D126", X"D12D", 
X"D134", X"D13B", X"D142", X"D149", X"D14F", X"D156", X"D15D", X"D164", X"D16B", X"D172", 
X"D179", X"D180", X"D187", X"D18D", X"D194", X"D19B", X"D1A2", X"D1A9", X"D1B0", X"D1B7", 
X"D1BE", X"D1C5", X"D1CB", X"D1D2", X"D1D9", X"D1E0", X"D1E7", X"D1EE", X"D1F5", X"D1FB", 
X"D202", X"D209", X"D210", X"D217", X"D21E", X"D225", X"D22B", X"D232", X"D239", X"D240", 
X"D247", X"D24E", X"D255", X"D25B", X"D262", X"D269", X"D270", X"D277", X"D27E", X"D284", 
X"D28B", X"D292", X"D299", X"D2A0", X"D2A7", X"D2AD", X"D2B4", X"D2BB", X"D2C2", X"D2C9", 
X"D2CF", X"D2D6", X"D2DD", X"D2E4", X"D2EB", X"D2F2", X"D2F8", X"D2FF", X"D306", X"D30D", 
X"D314", X"D31A", X"D321", X"D328", X"D32F", X"D335", X"D33C", X"D343", X"D34A", X"D351", 
X"D357", X"D35E", X"D365", X"D36C", X"D373", X"D379", X"D380", X"D387", X"D38E", X"D394", 
X"D39B", X"D3A2", X"D3A9", X"D3AF", X"D3B6", X"D3BD", X"D3C4", X"D3CA", X"D3D1", X"D3D8", 
X"D3DF", X"D3E6", X"D3EC", X"D3F3", X"D3FA", X"D400", X"D407", X"D40E", X"D415", X"D41B", 
X"D422", X"D429", X"D430", X"D436", X"D43D", X"D444", X"D44B", X"D451", X"D458", X"D45F", 
X"D465", X"D46C", X"D473", X"D47A", X"D480", X"D487", X"D48E", X"D494", X"D49B", X"D4A2", 
X"D4A9", X"D4AF", X"D4B6", X"D4BD", X"D4C3", X"D4CA", X"D4D1", X"D4D7", X"D4DE", X"D4E5", 
X"D4EB", X"D4F2", X"D4F9", X"D500", X"D506", X"D50D", X"D514", X"D51A", X"D521", X"D528", 
X"D52E", X"D535", X"D53C", X"D542", X"D549", X"D550", X"D556", X"D55D", X"D564", X"D56A", 
X"D571", X"D578", X"D57E", X"D585", X"D58B", X"D592", X"D599", X"D59F", X"D5A6", X"D5AD", 
X"D5B3", X"D5BA", X"D5C1", X"D5C7", X"D5CE", X"D5D5", X"D5DB", X"D5E2", X"D5E8", X"D5EF", 
X"D5F6", X"D5FC", X"D603", X"D60A", X"D610", X"D617", X"D61D", X"D624", X"D62B", X"D631", 
X"D638", X"D63E", X"D645", X"D64C", X"D652", X"D659", X"D65F", X"D666", X"D66D", X"D673", 
X"D67A", X"D680", X"D687", X"D68D", X"D694", X"D69B", X"D6A1", X"D6A8", X"D6AE", X"D6B5", 
X"D6BC", X"D6C2", X"D6C9", X"D6CF", X"D6D6", X"D6DC", X"D6E3", X"D6EA", X"D6F0", X"D6F7", 
X"D6FD", X"D704", X"D70A", X"D711", X"D717", X"D71E", X"D724", X"D72B", X"D732", X"D738", 
X"D73F", X"D745", X"D74C", X"D752", X"D759", X"D75F", X"D766", X"D76C", X"D773", X"D779", 
X"D780", X"D786", X"D78D", X"D794", X"D79A", X"D7A1", X"D7A7", X"D7AE", X"D7B4", X"D7BB", 
X"D7C1", X"D7C8", X"D7CE", X"D7D5", X"D7DB", X"D7E2", X"D7E8", X"D7EF", X"D7F5", X"D7FC", 
X"D802", X"D809", X"D80F", X"D816", X"D81C", X"D822", X"D829", X"D82F", X"D836", X"D83C", 
X"D843", X"D849", X"D850", X"D856", X"D85D", X"D863", X"D86A", X"D870", X"D877", X"D87D", 
X"D884", X"D88A", X"D890", X"D897", X"D89D", X"D8A4", X"D8AA", X"D8B1", X"D8B7", X"D8BE", 
X"D8C4", X"D8CA", X"D8D1", X"D8D7", X"D8DE", X"D8E4", X"D8EB", X"D8F1", X"D8F7", X"D8FE", 
X"D904", X"D90B", X"D911", X"D918", X"D91E", X"D924", X"D92B", X"D931", X"D938", X"D93E", 
X"D944", X"D94B", X"D951", X"D958", X"D95E", X"D964", X"D96B", X"D971", X"D978", X"D97E", 
X"D984", X"D98B", X"D991", X"D998", X"D99E", X"D9A4", X"D9AB", X"D9B1", X"D9B7", X"D9BE", 
X"D9C4", X"D9CB", X"D9D1", X"D9D7", X"D9DE", X"D9E4", X"D9EA", X"D9F1", X"D9F7", X"D9FD", 
X"DA04", X"DA0A", X"DA10", X"DA17", X"DA1D", X"DA24", X"DA2A", X"DA30", X"DA37", X"DA3D", 
X"DA43", X"DA4A", X"DA50", X"DA56", X"DA5D", X"DA63", X"DA69", X"DA70", X"DA76", X"DA7C", 
X"DA82", X"DA89", X"DA8F", X"DA95", X"DA9C", X"DAA2", X"DAA8", X"DAAF", X"DAB5", X"DABB", 
X"DAC2", X"DAC8", X"DACE", X"DAD4", X"DADB", X"DAE1", X"DAE7", X"DAEE", X"DAF4", X"DAFA", 
X"DB01", X"DB07", X"DB0D", X"DB13", X"DB1A", X"DB20", X"DB26", X"DB2C", X"DB33", X"DB39", 
X"DB3F", X"DB46", X"DB4C", X"DB52", X"DB58", X"DB5F", X"DB65", X"DB6B", X"DB71", X"DB78", 
X"DB7E", X"DB84", X"DB8A", X"DB91", X"DB97", X"DB9D", X"DBA3", X"DBAA", X"DBB0", X"DBB6", 
X"DBBC", X"DBC2", X"DBC9", X"DBCF", X"DBD5", X"DBDB", X"DBE2", X"DBE8", X"DBEE", X"DBF4", 
X"DBFA", X"DC01", X"DC07", X"DC0D", X"DC13", X"DC1A", X"DC20", X"DC26", X"DC2C", X"DC32", 
X"DC39", X"DC3F", X"DC45", X"DC4B", X"DC51", X"DC58", X"DC5E", X"DC64", X"DC6A", X"DC70", 
X"DC76", X"DC7D", X"DC83", X"DC89", X"DC8F", X"DC95", X"DC9B", X"DCA2", X"DCA8", X"DCAE", 
X"DCB4", X"DCBA", X"DCC0", X"DCC7", X"DCCD", X"DCD3", X"DCD9", X"DCDF", X"DCE5", X"DCEC", 
X"DCF2", X"DCF8", X"DCFE", X"DD04", X"DD0A", X"DD10", X"DD16", X"DD1D", X"DD23", X"DD29", 
X"DD2F", X"DD35", X"DD3B", X"DD41", X"DD48", X"DD4E", X"DD54", X"DD5A", X"DD60", X"DD66", 
X"DD6C", X"DD72", X"DD78", X"DD7F", X"DD85", X"DD8B", X"DD91", X"DD97", X"DD9D", X"DDA3", 
X"DDA9", X"DDAF", X"DDB5", X"DDBB", X"DDC2", X"DDC8", X"DDCE", X"DDD4", X"DDDA", X"DDE0", 
X"DDE6", X"DDEC", X"DDF2", X"DDF8", X"DDFE", X"DE04", X"DE0A", X"DE10", X"DE17", X"DE1D", 
X"DE23", X"DE29", X"DE2F", X"DE35", X"DE3B", X"DE41", X"DE47", X"DE4D", X"DE53", X"DE59", 
X"DE5F", X"DE65", X"DE6B", X"DE71", X"DE77", X"DE7D", X"DE83", X"DE89", X"DE8F", X"DE95", 
X"DE9B", X"DEA1", X"DEA7", X"DEAD", X"DEB3", X"DEB9", X"DEBF", X"DEC5", X"DECB", X"DED1", 
X"DED7", X"DEDD", X"DEE3", X"DEE9", X"DEEF", X"DEF5", X"DEFB", X"DF01", X"DF07", X"DF0D", 
X"DF13", X"DF19", X"DF1F", X"DF25", X"DF2B", X"DF31", X"DF37", X"DF3D", X"DF43", X"DF49", 
X"DF4F", X"DF55", X"DF5B", X"DF61", X"DF67", X"DF6D", X"DF73", X"DF79", X"DF7F", X"DF85", 
X"DF8B", X"DF91", X"DF97", X"DF9D", X"DFA2", X"DFA8", X"DFAE", X"DFB4", X"DFBA", X"DFC0", 
X"DFC6", X"DFCC", X"DFD2", X"DFD8", X"DFDE", X"DFE4", X"DFEA", X"DFF0", X"DFF5", X"DFFB", 
X"E001", X"E007", X"E00D", X"E013", X"E019", X"E01F", X"E025", X"E02B", X"E031", X"E036", 
X"E03C", X"E042", X"E048", X"E04E", X"E054", X"E05A", X"E060", X"E065", X"E06B", X"E071", 
X"E077", X"E07D", X"E083", X"E089", X"E08F", X"E094", X"E09A", X"E0A0", X"E0A6", X"E0AC", 
X"E0B2", X"E0B8", X"E0BD", X"E0C3", X"E0C9", X"E0CF", X"E0D5", X"E0DB", X"E0E1", X"E0E6", 
X"E0EC", X"E0F2", X"E0F8", X"E0FE", X"E104", X"E109", X"E10F", X"E115", X"E11B", X"E121", 
X"E126", X"E12C", X"E132", X"E138", X"E13E", X"E144", X"E149", X"E14F", X"E155", X"E15B", 
X"E161", X"E166", X"E16C", X"E172", X"E178", X"E17E", X"E183", X"E189", X"E18F", X"E195", 
X"E19A", X"E1A0", X"E1A6", X"E1AC", X"E1B2", X"E1B7", X"E1BD", X"E1C3", X"E1C9", X"E1CE", 
X"E1D4", X"E1DA", X"E1E0", X"E1E5", X"E1EB", X"E1F1", X"E1F7", X"E1FD", X"E202", X"E208", 
X"E20E", X"E213", X"E219", X"E21F", X"E225", X"E22A", X"E230", X"E236", X"E23C", X"E241", 
X"E247", X"E24D", X"E253", X"E258", X"E25E", X"E264", X"E269", X"E26F", X"E275", X"E27B", 
X"E280", X"E286", X"E28C", X"E291", X"E297", X"E29D", X"E2A2", X"E2A8", X"E2AE", X"E2B4", 
X"E2B9", X"E2BF", X"E2C5", X"E2CA", X"E2D0", X"E2D6", X"E2DB", X"E2E1", X"E2E7", X"E2EC", 
X"E2F2", X"E2F8", X"E2FD", X"E303", X"E309", X"E30E", X"E314", X"E31A", X"E31F", X"E325", 
X"E32B", X"E330", X"E336", X"E33C", X"E341", X"E347", X"E34C", X"E352", X"E358", X"E35D", 
X"E363", X"E369", X"E36E", X"E374", X"E37A", X"E37F", X"E385", X"E38A", X"E390", X"E396", 
X"E39B", X"E3A1", X"E3A6", X"E3AC", X"E3B2", X"E3B7", X"E3BD", X"E3C2", X"E3C8", X"E3CE", 
X"E3D3", X"E3D9", X"E3DE", X"E3E4", X"E3EA", X"E3EF", X"E3F5", X"E3FA", X"E400", X"E406", 
X"E40B", X"E411", X"E416", X"E41C", X"E421", X"E427", X"E42D", X"E432", X"E438", X"E43D", 
X"E443", X"E448", X"E44E", X"E453", X"E459", X"E45E", X"E464", X"E46A", X"E46F", X"E475", 
X"E47A", X"E480", X"E485", X"E48B", X"E490", X"E496", X"E49B", X"E4A1", X"E4A6", X"E4AC", 
X"E4B1", X"E4B7", X"E4BC", X"E4C2", X"E4C8", X"E4CD", X"E4D3", X"E4D8", X"E4DE", X"E4E3", 
X"E4E9", X"E4EE", X"E4F4", X"E4F9", X"E4FF", X"E504", X"E509", X"E50F", X"E514", X"E51A", 
X"E51F", X"E525", X"E52A", X"E530", X"E535", X"E53B", X"E540", X"E546", X"E54B", X"E551", 
X"E556", X"E55C", X"E561", X"E566", X"E56C", X"E571", X"E577", X"E57C", X"E582", X"E587", 
X"E58D", X"E592", X"E597", X"E59D", X"E5A2", X"E5A8", X"E5AD", X"E5B3", X"E5B8", X"E5BD", 
X"E5C3", X"E5C8", X"E5CE", X"E5D3", X"E5D9", X"E5DE", X"E5E3", X"E5E9", X"E5EE", X"E5F4", 
X"E5F9", X"E5FE", X"E604", X"E609", X"E60F", X"E614", X"E619", X"E61F", X"E624", X"E62A", 
X"E62F", X"E634", X"E63A", X"E63F", X"E644", X"E64A", X"E64F", X"E655", X"E65A", X"E65F", 
X"E665", X"E66A", X"E66F", X"E675", X"E67A", X"E67F", X"E685", X"E68A", X"E68F", X"E695", 
X"E69A", X"E6A0", X"E6A5", X"E6AA", X"E6B0", X"E6B5", X"E6BA", X"E6C0", X"E6C5", X"E6CA", 
X"E6D0", X"E6D5", X"E6DA", X"E6DF", X"E6E5", X"E6EA", X"E6EF", X"E6F5", X"E6FA", X"E6FF", 
X"E705", X"E70A", X"E70F", X"E715", X"E71A", X"E71F", X"E724", X"E72A", X"E72F", X"E734", 
X"E73A", X"E73F", X"E744", X"E749", X"E74F", X"E754", X"E759", X"E75F", X"E764", X"E769", 
X"E76E", X"E774", X"E779", X"E77E", X"E783", X"E789", X"E78E", X"E793", X"E798", X"E79E", 
X"E7A3", X"E7A8", X"E7AD", X"E7B3", X"E7B8", X"E7BD", X"E7C2", X"E7C8", X"E7CD", X"E7D2", 
X"E7D7", X"E7DC", X"E7E2", X"E7E7", X"E7EC", X"E7F1", X"E7F7", X"E7FC", X"E801", X"E806", 
X"E80B", X"E811", X"E816", X"E81B", X"E820", X"E825", X"E82B", X"E830", X"E835", X"E83A", 
X"E83F", X"E844", X"E84A", X"E84F", X"E854", X"E859", X"E85E", X"E864", X"E869", X"E86E", 
X"E873", X"E878", X"E87D", X"E883", X"E888", X"E88D", X"E892", X"E897", X"E89C", X"E8A1", 
X"E8A7", X"E8AC", X"E8B1", X"E8B6", X"E8BB", X"E8C0", X"E8C5", X"E8CB", X"E8D0", X"E8D5", 
X"E8DA", X"E8DF", X"E8E4", X"E8E9", X"E8EE", X"E8F4", X"E8F9", X"E8FE", X"E903", X"E908", 
X"E90D", X"E912", X"E917", X"E91C", X"E922", X"E927", X"E92C", X"E931", X"E936", X"E93B", 
X"E940", X"E945", X"E94A", X"E94F", X"E954", X"E959", X"E95F", X"E964", X"E969", X"E96E", 
X"E973", X"E978", X"E97D", X"E982", X"E987", X"E98C", X"E991", X"E996", X"E99B", X"E9A0", 
X"E9A5", X"E9AA", X"E9AF", X"E9B5", X"E9BA", X"E9BF", X"E9C4", X"E9C9", X"E9CE", X"E9D3", 
X"E9D8", X"E9DD", X"E9E2", X"E9E7", X"E9EC", X"E9F1", X"E9F6", X"E9FB", X"EA00", X"EA05", 
X"EA0A", X"EA0F", X"EA14", X"EA19", X"EA1E", X"EA23", X"EA28", X"EA2D", X"EA32", X"EA37", 
X"EA3C", X"EA41", X"EA46", X"EA4B", X"EA50", X"EA55", X"EA5A", X"EA5F", X"EA64", X"EA69", 
X"EA6E", X"EA73", X"EA78", X"EA7C", X"EA81", X"EA86", X"EA8B", X"EA90", X"EA95", X"EA9A", 
X"EA9F", X"EAA4", X"EAA9", X"EAAE", X"EAB3", X"EAB8", X"EABD", X"EAC2", X"EAC7", X"EACC", 
X"EAD0", X"EAD5", X"EADA", X"EADF", X"EAE4", X"EAE9", X"EAEE", X"EAF3", X"EAF8", X"EAFD", 
X"EB02", X"EB07", X"EB0B", X"EB10", X"EB15", X"EB1A", X"EB1F", X"EB24", X"EB29", X"EB2E", 
X"EB33", X"EB37", X"EB3C", X"EB41", X"EB46", X"EB4B", X"EB50", X"EB55", X"EB5A", X"EB5E", 
X"EB63", X"EB68", X"EB6D", X"EB72", X"EB77", X"EB7C", X"EB80", X"EB85", X"EB8A", X"EB8F", 
X"EB94", X"EB99", X"EB9D", X"EBA2", X"EBA7", X"EBAC", X"EBB1", X"EBB6", X"EBBA", X"EBBF", 
X"EBC4", X"EBC9", X"EBCE", X"EBD3", X"EBD7", X"EBDC", X"EBE1", X"EBE6", X"EBEB", X"EBEF", 
X"EBF4", X"EBF9", X"EBFE", X"EC03", X"EC07", X"EC0C", X"EC11", X"EC16", X"EC1B", X"EC1F", 
X"EC24", X"EC29", X"EC2E", X"EC32", X"EC37", X"EC3C", X"EC41", X"EC46", X"EC4A", X"EC4F", 
X"EC54", X"EC59", X"EC5D", X"EC62", X"EC67", X"EC6C", X"EC70", X"EC75", X"EC7A", X"EC7F", 
X"EC83", X"EC88", X"EC8D", X"EC92", X"EC96", X"EC9B", X"ECA0", X"ECA4", X"ECA9", X"ECAE", 
X"ECB3", X"ECB7", X"ECBC", X"ECC1", X"ECC6", X"ECCA", X"ECCF", X"ECD4", X"ECD8", X"ECDD", 
X"ECE2", X"ECE6", X"ECEB", X"ECF0", X"ECF5", X"ECF9", X"ECFE", X"ED03", X"ED07", X"ED0C", 
X"ED11", X"ED15", X"ED1A", X"ED1F", X"ED23", X"ED28", X"ED2D", X"ED31", X"ED36", X"ED3B", 
X"ED3F", X"ED44", X"ED49", X"ED4D", X"ED52", X"ED57", X"ED5B", X"ED60", X"ED64", X"ED69", 
X"ED6E", X"ED72", X"ED77", X"ED7C", X"ED80", X"ED85", X"ED8A", X"ED8E", X"ED93", X"ED97", 
X"ED9C", X"EDA1", X"EDA5", X"EDAA", X"EDAE", X"EDB3", X"EDB8", X"EDBC", X"EDC1", X"EDC5", 
X"EDCA", X"EDCF", X"EDD3", X"EDD8", X"EDDC", X"EDE1", X"EDE6", X"EDEA", X"EDEF", X"EDF3", 
X"EDF8", X"EDFC", X"EE01", X"EE06", X"EE0A", X"EE0F", X"EE13", X"EE18", X"EE1C", X"EE21", 
X"EE26", X"EE2A", X"EE2F", X"EE33", X"EE38", X"EE3C", X"EE41", X"EE45", X"EE4A", X"EE4E", 
X"EE53", X"EE57", X"EE5C", X"EE61", X"EE65", X"EE6A", X"EE6E", X"EE73", X"EE77", X"EE7C", 
X"EE80", X"EE85", X"EE89", X"EE8E", X"EE92", X"EE97", X"EE9B", X"EEA0", X"EEA4", X"EEA9", 
X"EEAD", X"EEB2", X"EEB6", X"EEBB", X"EEBF", X"EEC4", X"EEC8", X"EECD", X"EED1", X"EED5", 
X"EEDA", X"EEDE", X"EEE3", X"EEE7", X"EEEC", X"EEF0", X"EEF5", X"EEF9", X"EEFE", X"EF02", 
X"EF06", X"EF0B", X"EF0F", X"EF14", X"EF18", X"EF1D", X"EF21", X"EF26", X"EF2A", X"EF2E", 
X"EF33", X"EF37", X"EF3C", X"EF40", X"EF45", X"EF49", X"EF4D", X"EF52", X"EF56", X"EF5B", 
X"EF5F", X"EF63", X"EF68", X"EF6C", X"EF71", X"EF75", X"EF79", X"EF7E", X"EF82", X"EF87", 
X"EF8B", X"EF8F", X"EF94", X"EF98", X"EF9C", X"EFA1", X"EFA5", X"EFAA", X"EFAE", X"EFB2", 
X"EFB7", X"EFBB", X"EFBF", X"EFC4", X"EFC8", X"EFCC", X"EFD1", X"EFD5", X"EFDA", X"EFDE", 
X"EFE2", X"EFE7", X"EFEB", X"EFEF", X"EFF4", X"EFF8", X"EFFC", X"F001", X"F005", X"F009", 
X"F00D", X"F012", X"F016", X"F01A", X"F01F", X"F023", X"F027", X"F02C", X"F030", X"F034", 
X"F039", X"F03D", X"F041", X"F045", X"F04A", X"F04E", X"F052", X"F057", X"F05B", X"F05F", 
X"F063", X"F068", X"F06C", X"F070", X"F075", X"F079", X"F07D", X"F081", X"F086", X"F08A", 
X"F08E", X"F092", X"F097", X"F09B", X"F09F", X"F0A3", X"F0A8", X"F0AC", X"F0B0", X"F0B4", 
X"F0B9", X"F0BD", X"F0C1", X"F0C5", X"F0C9", X"F0CE", X"F0D2", X"F0D6", X"F0DA", X"F0DF", 
X"F0E3", X"F0E7", X"F0EB", X"F0EF", X"F0F4", X"F0F8", X"F0FC", X"F100", X"F104", X"F109", 
X"F10D", X"F111", X"F115", X"F119", X"F11E", X"F122", X"F126", X"F12A", X"F12E", X"F132", 
X"F137", X"F13B", X"F13F", X"F143", X"F147", X"F14B", X"F150", X"F154", X"F158", X"F15C", 
X"F160", X"F164", X"F168", X"F16D", X"F171", X"F175", X"F179", X"F17D", X"F181", X"F185", 
X"F18A", X"F18E", X"F192", X"F196", X"F19A", X"F19E", X"F1A2", X"F1A6", X"F1AB", X"F1AF", 
X"F1B3", X"F1B7", X"F1BB", X"F1BF", X"F1C3", X"F1C7", X"F1CB", X"F1CF", X"F1D3", X"F1D8", 
X"F1DC", X"F1E0", X"F1E4", X"F1E8", X"F1EC", X"F1F0", X"F1F4", X"F1F8", X"F1FC", X"F200", 
X"F204", X"F208", X"F20D", X"F211", X"F215", X"F219", X"F21D", X"F221", X"F225", X"F229", 
X"F22D", X"F231", X"F235", X"F239", X"F23D", X"F241", X"F245", X"F249", X"F24D", X"F251", 
X"F255", X"F259", X"F25D", X"F261", X"F265", X"F269", X"F26D", X"F271", X"F275", X"F279", 
X"F27D", X"F281", X"F285", X"F289", X"F28D", X"F291", X"F295", X"F299", X"F29D", X"F2A1", 
X"F2A5", X"F2A9", X"F2AD", X"F2B1", X"F2B5", X"F2B9", X"F2BD", X"F2C1", X"F2C5", X"F2C9", 
X"F2CD", X"F2D1", X"F2D5", X"F2D9", X"F2DD", X"F2E0", X"F2E4", X"F2E8", X"F2EC", X"F2F0", 
X"F2F4", X"F2F8", X"F2FC", X"F300", X"F304", X"F308", X"F30C", X"F310", X"F314", X"F317", 
X"F31B", X"F31F", X"F323", X"F327", X"F32B", X"F32F", X"F333", X"F337", X"F33B", X"F33E", 
X"F342", X"F346", X"F34A", X"F34E", X"F352", X"F356", X"F35A", X"F35D", X"F361", X"F365", 
X"F369", X"F36D", X"F371", X"F375", X"F379", X"F37C", X"F380", X"F384", X"F388", X"F38C", 
X"F390", X"F393", X"F397", X"F39B", X"F39F", X"F3A3", X"F3A7", X"F3AA", X"F3AE", X"F3B2", 
X"F3B6", X"F3BA", X"F3BE", X"F3C1", X"F3C5", X"F3C9", X"F3CD", X"F3D1", X"F3D4", X"F3D8", 
X"F3DC", X"F3E0", X"F3E4", X"F3E7", X"F3EB", X"F3EF", X"F3F3", X"F3F7", X"F3FA", X"F3FE", 
X"F402", X"F406", X"F409", X"F40D", X"F411", X"F415", X"F419", X"F41C", X"F420", X"F424", 
X"F428", X"F42B", X"F42F", X"F433", X"F437", X"F43A", X"F43E", X"F442", X"F446", X"F449", 
X"F44D", X"F451", X"F454", X"F458", X"F45C", X"F460", X"F463", X"F467", X"F46B", X"F46E", 
X"F472", X"F476", X"F47A", X"F47D", X"F481", X"F485", X"F488", X"F48C", X"F490", X"F493", 
X"F497", X"F49B", X"F49F", X"F4A2", X"F4A6", X"F4AA", X"F4AD", X"F4B1", X"F4B5", X"F4B8", 
X"F4BC", X"F4C0", X"F4C3", X"F4C7", X"F4CB", X"F4CE", X"F4D2", X"F4D6", X"F4D9", X"F4DD", 
X"F4E1", X"F4E4", X"F4E8", X"F4EB", X"F4EF", X"F4F3", X"F4F6", X"F4FA", X"F4FE", X"F501", 
X"F505", X"F508", X"F50C", X"F510", X"F513", X"F517", X"F51B", X"F51E", X"F522", X"F525", 
X"F529", X"F52D", X"F530", X"F534", X"F537", X"F53B", X"F53E", X"F542", X"F546", X"F549", 
X"F54D", X"F550", X"F554", X"F558", X"F55B", X"F55F", X"F562", X"F566", X"F569", X"F56D", 
X"F570", X"F574", X"F578", X"F57B", X"F57F", X"F582", X"F586", X"F589", X"F58D", X"F590", 
X"F594", X"F597", X"F59B", X"F59E", X"F5A2", X"F5A6", X"F5A9", X"F5AD", X"F5B0", X"F5B4", 
X"F5B7", X"F5BB", X"F5BE", X"F5C2", X"F5C5", X"F5C9", X"F5CC", X"F5D0", X"F5D3", X"F5D7", 
X"F5DA", X"F5DE", X"F5E1", X"F5E5", X"F5E8", X"F5EB", X"F5EF", X"F5F2", X"F5F6", X"F5F9", 
X"F5FD", X"F600", X"F604", X"F607", X"F60B", X"F60E", X"F612", X"F615", X"F618", X"F61C", 
X"F61F", X"F623", X"F626", X"F62A", X"F62D", X"F631", X"F634", X"F637", X"F63B", X"F63E", 
X"F642", X"F645", X"F649", X"F64C", X"F64F", X"F653", X"F656", X"F65A", X"F65D", X"F660", 
X"F664", X"F667", X"F66B", X"F66E", X"F671", X"F675", X"F678", X"F67B", X"F67F", X"F682", 
X"F686", X"F689", X"F68C", X"F690", X"F693", X"F696", X"F69A", X"F69D", X"F6A1", X"F6A4", 
X"F6A7", X"F6AB", X"F6AE", X"F6B1", X"F6B5", X"F6B8", X"F6BB", X"F6BF", X"F6C2", X"F6C5", 
X"F6C9", X"F6CC", X"F6CF", X"F6D3", X"F6D6", X"F6D9", X"F6DD", X"F6E0", X"F6E3", X"F6E7", 
X"F6EA", X"F6ED", X"F6F0", X"F6F4", X"F6F7", X"F6FA", X"F6FE", X"F701", X"F704", X"F708", 
X"F70B", X"F70E", X"F711", X"F715", X"F718", X"F71B", X"F71E", X"F722", X"F725", X"F728", 
X"F72C", X"F72F", X"F732", X"F735", X"F739", X"F73C", X"F73F", X"F742", X"F746", X"F749", 
X"F74C", X"F74F", X"F753", X"F756", X"F759", X"F75C", X"F75F", X"F763", X"F766", X"F769", 
X"F76C", X"F770", X"F773", X"F776", X"F779", X"F77C", X"F780", X"F783", X"F786", X"F789", 
X"F78C", X"F790", X"F793", X"F796", X"F799", X"F79C", X"F79F", X"F7A3", X"F7A6", X"F7A9", 
X"F7AC", X"F7AF", X"F7B3", X"F7B6", X"F7B9", X"F7BC", X"F7BF", X"F7C2", X"F7C5", X"F7C9", 
X"F7CC", X"F7CF", X"F7D2", X"F7D5", X"F7D8", X"F7DB", X"F7DF", X"F7E2", X"F7E5", X"F7E8", 
X"F7EB", X"F7EE", X"F7F1", X"F7F4", X"F7F8", X"F7FB", X"F7FE", X"F801", X"F804", X"F807", 
X"F80A", X"F80D", X"F810", X"F814", X"F817", X"F81A", X"F81D", X"F820", X"F823", X"F826", 
X"F829", X"F82C", X"F82F", X"F832", X"F835", X"F839", X"F83C", X"F83F", X"F842", X"F845", 
X"F848", X"F84B", X"F84E", X"F851", X"F854", X"F857", X"F85A", X"F85D", X"F860", X"F863", 
X"F866", X"F869", X"F86C", X"F86F", X"F872", X"F875", X"F878", X"F87B", X"F87E", X"F882", 
X"F885", X"F888", X"F88B", X"F88E", X"F891", X"F894", X"F897", X"F89A", X"F89D", X"F8A0", 
X"F8A3", X"F8A5", X"F8A8", X"F8AB", X"F8AE", X"F8B1", X"F8B4", X"F8B7", X"F8BA", X"F8BD", 
X"F8C0", X"F8C3", X"F8C6", X"F8C9", X"F8CC", X"F8CF", X"F8D2", X"F8D5", X"F8D8", X"F8DB", 
X"F8DE", X"F8E1", X"F8E4", X"F8E7", X"F8EA", X"F8EC", X"F8EF", X"F8F2", X"F8F5", X"F8F8", 
X"F8FB", X"F8FE", X"F901", X"F904", X"F907", X"F90A", X"F90D", X"F90F", X"F912", X"F915", 
X"F918", X"F91B", X"F91E", X"F921", X"F924", X"F927", X"F929", X"F92C", X"F92F", X"F932", 
X"F935", X"F938", X"F93B", X"F93E", X"F940", X"F943", X"F946", X"F949", X"F94C", X"F94F", 
X"F952", X"F954", X"F957", X"F95A", X"F95D", X"F960", X"F963", X"F966", X"F968", X"F96B", 
X"F96E", X"F971", X"F974", X"F976", X"F979", X"F97C", X"F97F", X"F982", X"F985", X"F987", 
X"F98A", X"F98D", X"F990", X"F993", X"F995", X"F998", X"F99B", X"F99E", X"F9A0", X"F9A3", 
X"F9A6", X"F9A9", X"F9AC", X"F9AE", X"F9B1", X"F9B4", X"F9B7", X"F9B9", X"F9BC", X"F9BF", 
X"F9C2", X"F9C4", X"F9C7", X"F9CA", X"F9CD", X"F9CF", X"F9D2", X"F9D5", X"F9D8", X"F9DA", 
X"F9DD", X"F9E0", X"F9E3", X"F9E5", X"F9E8", X"F9EB", X"F9EE", X"F9F0", X"F9F3", X"F9F6", 
X"F9F8", X"F9FB", X"F9FE", X"FA01", X"FA03", X"FA06", X"FA09", X"FA0B", X"FA0E", X"FA11", 
X"FA13", X"FA16", X"FA19", X"FA1B", X"FA1E", X"FA21", X"FA23", X"FA26", X"FA29", X"FA2B", 
X"FA2E", X"FA31", X"FA33", X"FA36", X"FA39", X"FA3B", X"FA3E", X"FA41", X"FA43", X"FA46", 
X"FA49", X"FA4B", X"FA4E", X"FA51", X"FA53", X"FA56", X"FA58", X"FA5B", X"FA5E", X"FA60", 
X"FA63", X"FA66", X"FA68", X"FA6B", X"FA6D", X"FA70", X"FA73", X"FA75", X"FA78", X"FA7A", 
X"FA7D", X"FA80", X"FA82", X"FA85", X"FA87", X"FA8A", X"FA8D", X"FA8F", X"FA92", X"FA94", 
X"FA97", X"FA99", X"FA9C", X"FA9F", X"FAA1", X"FAA4", X"FAA6", X"FAA9", X"FAAB", X"FAAE", 
X"FAB0", X"FAB3", X"FAB6", X"FAB8", X"FABB", X"FABD", X"FAC0", X"FAC2", X"FAC5", X"FAC7", 
X"FACA", X"FACC", X"FACF", X"FAD1", X"FAD4", X"FAD6", X"FAD9", X"FADB", X"FADE", X"FAE0", 
X"FAE3", X"FAE5", X"FAE8", X"FAEA", X"FAED", X"FAEF", X"FAF2", X"FAF4", X"FAF7", X"FAF9", 
X"FAFC", X"FAFE", X"FB01", X"FB03", X"FB06", X"FB08", X"FB0B", X"FB0D", X"FB10", X"FB12", 
X"FB14", X"FB17", X"FB19", X"FB1C", X"FB1E", X"FB21", X"FB23", X"FB26", X"FB28", X"FB2A", 
X"FB2D", X"FB2F", X"FB32", X"FB34", X"FB37", X"FB39", X"FB3B", X"FB3E", X"FB40", X"FB43", 
X"FB45", X"FB47", X"FB4A", X"FB4C", X"FB4F", X"FB51", X"FB53", X"FB56", X"FB58", X"FB5B", 
X"FB5D", X"FB5F", X"FB62", X"FB64", X"FB67", X"FB69", X"FB6B", X"FB6E", X"FB70", X"FB72", 
X"FB75", X"FB77", X"FB79", X"FB7C", X"FB7E", X"FB81", X"FB83", X"FB85", X"FB88", X"FB8A", 
X"FB8C", X"FB8F", X"FB91", X"FB93", X"FB96", X"FB98", X"FB9A", X"FB9D", X"FB9F", X"FBA1", 
X"FBA3", X"FBA6", X"FBA8", X"FBAA", X"FBAD", X"FBAF", X"FBB1", X"FBB4", X"FBB6", X"FBB8", 
X"FBBA", X"FBBD", X"FBBF", X"FBC1", X"FBC4", X"FBC6", X"FBC8", X"FBCA", X"FBCD", X"FBCF", 
X"FBD1", X"FBD4", X"FBD6", X"FBD8", X"FBDA", X"FBDD", X"FBDF", X"FBE1", X"FBE3", X"FBE6", 
X"FBE8", X"FBEA", X"FBEC", X"FBEE", X"FBF1", X"FBF3", X"FBF5", X"FBF7", X"FBFA", X"FBFC", 
X"FBFE", X"FC00", X"FC03", X"FC05", X"FC07", X"FC09", X"FC0B", X"FC0E", X"FC10", X"FC12", 
X"FC14", X"FC16", X"FC19", X"FC1B", X"FC1D", X"FC1F", X"FC21", X"FC23", X"FC26", X"FC28", 
X"FC2A", X"FC2C", X"FC2E", X"FC30", X"FC33", X"FC35", X"FC37", X"FC39", X"FC3B", X"FC3D", 
X"FC40", X"FC42", X"FC44", X"FC46", X"FC48", X"FC4A", X"FC4C", X"FC4F", X"FC51", X"FC53", 
X"FC55", X"FC57", X"FC59", X"FC5B", X"FC5D", X"FC60", X"FC62", X"FC64", X"FC66", X"FC68", 
X"FC6A", X"FC6C", X"FC6E", X"FC70", X"FC72", X"FC75", X"FC77", X"FC79", X"FC7B", X"FC7D", 
X"FC7F", X"FC81", X"FC83", X"FC85", X"FC87", X"FC89", X"FC8B", X"FC8D", X"FC8F", X"FC92", 
X"FC94", X"FC96", X"FC98", X"FC9A", X"FC9C", X"FC9E", X"FCA0", X"FCA2", X"FCA4", X"FCA6", 
X"FCA8", X"FCAA", X"FCAC", X"FCAE", X"FCB0", X"FCB2", X"FCB4", X"FCB6", X"FCB8", X"FCBA", 
X"FCBC", X"FCBE", X"FCC0", X"FCC2", X"FCC4", X"FCC6", X"FCC8", X"FCCA", X"FCCC", X"FCCE", 
X"FCD0", X"FCD2", X"FCD4", X"FCD6", X"FCD8", X"FCDA", X"FCDC", X"FCDE", X"FCE0", X"FCE2", 
X"FCE4", X"FCE6", X"FCE8", X"FCEA", X"FCEC", X"FCEE", X"FCF0", X"FCF1", X"FCF3", X"FCF5", 
X"FCF7", X"FCF9", X"FCFB", X"FCFD", X"FCFF", X"FD01", X"FD03", X"FD05", X"FD07", X"FD09", 
X"FD0A", X"FD0C", X"FD0E", X"FD10", X"FD12", X"FD14", X"FD16", X"FD18", X"FD1A", X"FD1C", 
X"FD1D", X"FD1F", X"FD21", X"FD23", X"FD25", X"FD27", X"FD29", X"FD2B", X"FD2C", X"FD2E", 
X"FD30", X"FD32", X"FD34", X"FD36", X"FD38", X"FD3A", X"FD3B", X"FD3D", X"FD3F", X"FD41", 
X"FD43", X"FD45", X"FD46", X"FD48", X"FD4A", X"FD4C", X"FD4E", X"FD50", X"FD51", X"FD53", 
X"FD55", X"FD57", X"FD59", X"FD5A", X"FD5C", X"FD5E", X"FD60", X"FD62", X"FD63", X"FD65", 
X"FD67", X"FD69", X"FD6B", X"FD6C", X"FD6E", X"FD70", X"FD72", X"FD74", X"FD75", X"FD77", 
X"FD79", X"FD7B", X"FD7C", X"FD7E", X"FD80", X"FD82", X"FD83", X"FD85", X"FD87", X"FD89", 
X"FD8A", X"FD8C", X"FD8E", X"FD90", X"FD91", X"FD93", X"FD95", X"FD97", X"FD98", X"FD9A", 
X"FD9C", X"FD9D", X"FD9F", X"FDA1", X"FDA3", X"FDA4", X"FDA6", X"FDA8", X"FDA9", X"FDAB", 
X"FDAD", X"FDAE", X"FDB0", X"FDB2", X"FDB4", X"FDB5", X"FDB7", X"FDB9", X"FDBA", X"FDBC", 
X"FDBE", X"FDBF", X"FDC1", X"FDC3", X"FDC4", X"FDC6", X"FDC8", X"FDC9", X"FDCB", X"FDCD", 
X"FDCE", X"FDD0", X"FDD1", X"FDD3", X"FDD5", X"FDD6", X"FDD8", X"FDDA", X"FDDB", X"FDDD", 
X"FDDF", X"FDE0", X"FDE2", X"FDE3", X"FDE5", X"FDE7", X"FDE8", X"FDEA", X"FDEB", X"FDED", 
X"FDEF", X"FDF0", X"FDF2", X"FDF3", X"FDF5", X"FDF7", X"FDF8", X"FDFA", X"FDFB", X"FDFD", 
X"FDFF", X"FE00", X"FE02", X"FE03", X"FE05", X"FE06", X"FE08", X"FE0A", X"FE0B", X"FE0D", 
X"FE0E", X"FE10", X"FE11", X"FE13", X"FE14", X"FE16", X"FE17", X"FE19", X"FE1B", X"FE1C", 
X"FE1E", X"FE1F", X"FE21", X"FE22", X"FE24", X"FE25", X"FE27", X"FE28", X"FE2A", X"FE2B", 
X"FE2D", X"FE2E", X"FE30", X"FE31", X"FE33", X"FE34", X"FE36", X"FE37", X"FE39", X"FE3A", 
X"FE3C", X"FE3D", X"FE3F", X"FE40", X"FE42", X"FE43", X"FE44", X"FE46", X"FE47", X"FE49", 
X"FE4A", X"FE4C", X"FE4D", X"FE4F", X"FE50", X"FE52", X"FE53", X"FE54", X"FE56", X"FE57", 
X"FE59", X"FE5A", X"FE5C", X"FE5D", X"FE5E", X"FE60", X"FE61", X"FE63", X"FE64", X"FE66", 
X"FE67", X"FE68", X"FE6A", X"FE6B", X"FE6D", X"FE6E", X"FE6F", X"FE71", X"FE72", X"FE74", 
X"FE75", X"FE76", X"FE78", X"FE79", X"FE7A", X"FE7C", X"FE7D", X"FE7F", X"FE80", X"FE81", 
X"FE83", X"FE84", X"FE85", X"FE87", X"FE88", X"FE89", X"FE8B", X"FE8C", X"FE8D", X"FE8F", 
X"FE90", X"FE91", X"FE93", X"FE94", X"FE95", X"FE97", X"FE98", X"FE99", X"FE9B", X"FE9C", 
X"FE9D", X"FE9F", X"FEA0", X"FEA1", X"FEA3", X"FEA4", X"FEA5", X"FEA6", X"FEA8", X"FEA9", 
X"FEAA", X"FEAC", X"FEAD", X"FEAE", X"FEAF", X"FEB1", X"FEB2", X"FEB3", X"FEB5", X"FEB6", 
X"FEB7", X"FEB8", X"FEBA", X"FEBB", X"FEBC", X"FEBD", X"FEBF", X"FEC0", X"FEC1", X"FEC2", 
X"FEC4", X"FEC5", X"FEC6", X"FEC7", X"FEC9", X"FECA", X"FECB", X"FECC", X"FECD", X"FECF", 
X"FED0", X"FED1", X"FED2", X"FED3", X"FED5", X"FED6", X"FED7", X"FED8", X"FED9", X"FEDB", 
X"FEDC", X"FEDD", X"FEDE", X"FEDF", X"FEE1", X"FEE2", X"FEE3", X"FEE4", X"FEE5", X"FEE6", 
X"FEE8", X"FEE9", X"FEEA", X"FEEB", X"FEEC", X"FEED", X"FEEF", X"FEF0", X"FEF1", X"FEF2", 
X"FEF3", X"FEF4", X"FEF5", X"FEF7", X"FEF8", X"FEF9", X"FEFA", X"FEFB", X"FEFC", X"FEFD", 
X"FEFF", X"FF00", X"FF01", X"FF02", X"FF03", X"FF04", X"FF05", X"FF06", X"FF07", X"FF08", 
X"FF0A", X"FF0B", X"FF0C", X"FF0D", X"FF0E", X"FF0F", X"FF10", X"FF11", X"FF12", X"FF13", 
X"FF14", X"FF15", X"FF17", X"FF18", X"FF19", X"FF1A", X"FF1B", X"FF1C", X"FF1D", X"FF1E", 
X"FF1F", X"FF20", X"FF21", X"FF22", X"FF23", X"FF24", X"FF25", X"FF26", X"FF27", X"FF28", 
X"FF29", X"FF2A", X"FF2B", X"FF2C", X"FF2D", X"FF2E", X"FF2F", X"FF30", X"FF31", X"FF32", 
X"FF33", X"FF34", X"FF35", X"FF36", X"FF37", X"FF38", X"FF39", X"FF3A", X"FF3B", X"FF3C", 
X"FF3D", X"FF3E", X"FF3F", X"FF40", X"FF41", X"FF42", X"FF43", X"FF44", X"FF45", X"FF46", 
X"FF47", X"FF48", X"FF49", X"FF4A", X"FF4B", X"FF4C", X"FF4C", X"FF4D", X"FF4E", X"FF4F", 
X"FF50", X"FF51", X"FF52", X"FF53", X"FF54", X"FF55", X"FF56", X"FF57", X"FF58", X"FF58", 
X"FF59", X"FF5A", X"FF5B", X"FF5C", X"FF5D", X"FF5E", X"FF5F", X"FF60", X"FF60", X"FF61", 
X"FF62", X"FF63", X"FF64", X"FF65", X"FF66", X"FF67", X"FF67", X"FF68", X"FF69", X"FF6A", 
X"FF6B", X"FF6C", X"FF6D", X"FF6D", X"FF6E", X"FF6F", X"FF70", X"FF71", X"FF72", X"FF72", 
X"FF73", X"FF74", X"FF75", X"FF76", X"FF77", X"FF77", X"FF78", X"FF79", X"FF7A", X"FF7B", 
X"FF7B", X"FF7C", X"FF7D", X"FF7E", X"FF7F", X"FF7F", X"FF80", X"FF81", X"FF82", X"FF83", 
X"FF83", X"FF84", X"FF85", X"FF86", X"FF86", X"FF87", X"FF88", X"FF89", X"FF89", X"FF8A", 
X"FF8B", X"FF8C", X"FF8C", X"FF8D", X"FF8E", X"FF8F", X"FF8F", X"FF90", X"FF91", X"FF92", 
X"FF92", X"FF93", X"FF94", X"FF95", X"FF95", X"FF96", X"FF97", X"FF97", X"FF98", X"FF99", 
X"FF9A", X"FF9A", X"FF9B", X"FF9C", X"FF9C", X"FF9D", X"FF9E", X"FF9E", X"FF9F", X"FFA0", 
X"FFA1", X"FFA1", X"FFA2", X"FFA3", X"FFA3", X"FFA4", X"FFA5", X"FFA5", X"FFA6", X"FFA7", 
X"FFA7", X"FFA8", X"FFA9", X"FFA9", X"FFAA", X"FFAA", X"FFAB", X"FFAC", X"FFAC", X"FFAD", 
X"FFAE", X"FFAE", X"FFAF", X"FFB0", X"FFB0", X"FFB1", X"FFB1", X"FFB2", X"FFB3", X"FFB3", 
X"FFB4", X"FFB4", X"FFB5", X"FFB6", X"FFB6", X"FFB7", X"FFB7", X"FFB8", X"FFB9", X"FFB9", 
X"FFBA", X"FFBA", X"FFBB", X"FFBC", X"FFBC", X"FFBD", X"FFBD", X"FFBE", X"FFBE", X"FFBF", 
X"FFC0", X"FFC0", X"FFC1", X"FFC1", X"FFC2", X"FFC2", X"FFC3", X"FFC3", X"FFC4", X"FFC5", 
X"FFC5", X"FFC6", X"FFC6", X"FFC7", X"FFC7", X"FFC8", X"FFC8", X"FFC9", X"FFC9", X"FFCA", 
X"FFCA", X"FFCB", X"FFCB", X"FFCC", X"FFCC", X"FFCD", X"FFCD", X"FFCE", X"FFCE", X"FFCF", 
X"FFCF", X"FFD0", X"FFD0", X"FFD1", X"FFD1", X"FFD2", X"FFD2", X"FFD3", X"FFD3", X"FFD4", 
X"FFD4", X"FFD4", X"FFD5", X"FFD5", X"FFD6", X"FFD6", X"FFD7", X"FFD7", X"FFD8", X"FFD8", 
X"FFD9", X"FFD9", X"FFD9", X"FFDA", X"FFDA", X"FFDB", X"FFDB", X"FFDC", X"FFDC", X"FFDC", 
X"FFDD", X"FFDD", X"FFDE", X"FFDE", X"FFDE", X"FFDF", X"FFDF", X"FFE0", X"FFE0", X"FFE0", 
X"FFE1", X"FFE1", X"FFE2", X"FFE2", X"FFE2", X"FFE3", X"FFE3", X"FFE3", X"FFE4", X"FFE4", 
X"FFE5", X"FFE5", X"FFE5", X"FFE6", X"FFE6", X"FFE6", X"FFE7", X"FFE7", X"FFE7", X"FFE8", 
X"FFE8", X"FFE8", X"FFE9", X"FFE9", X"FFE9", X"FFEA", X"FFEA", X"FFEA", X"FFEB", X"FFEB", 
X"FFEB", X"FFEC", X"FFEC", X"FFEC", X"FFED", X"FFED", X"FFED", X"FFEE", X"FFEE", X"FFEE", 
X"FFEE", X"FFEF", X"FFEF", X"FFEF", X"FFF0", X"FFF0", X"FFF0", X"FFF0", X"FFF1", X"FFF1", 
X"FFF1", X"FFF2", X"FFF2", X"FFF2", X"FFF2", X"FFF3", X"FFF3", X"FFF3", X"FFF3", X"FFF4", 
X"FFF4", X"FFF4", X"FFF4", X"FFF5", X"FFF5", X"FFF5", X"FFF5", X"FFF5", X"FFF6", X"FFF6", 
X"FFF6", X"FFF6", X"FFF7", X"FFF7", X"FFF7", X"FFF7", X"FFF7", X"FFF8", X"FFF8", X"FFF8", 
X"FFF8", X"FFF8", X"FFF9", X"FFF9", X"FFF9", X"FFF9", X"FFF9", X"FFFA", X"FFFA", X"FFFA", 
X"FFFA", X"FFFA", X"FFFA", X"FFFB", X"FFFB", X"FFFB", X"FFFB", X"FFFB", X"FFFB", X"FFFB", 
X"FFFC", X"FFFC", X"FFFC", X"FFFC", X"FFFC", X"FFFC", X"FFFC", X"FFFD", X"FFFD", X"FFFD", 
X"FFFD", X"FFFD", X"FFFD", X"FFFD", X"FFFD", X"FFFE", X"FFFE", X"FFFE", X"FFFE", X"FFFE", 
X"FFFE", X"FFFE", X"FFFE", X"FFFE", X"FFFE", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", 
X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", 
X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", 
X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", 
X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", 
X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", 
X"8000", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", 
X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFF", X"FFFE", X"FFFE", X"FFFE", X"FFFE", 
X"FFFE", X"FFFE", X"FFFE", X"FFFE", X"FFFE", X"FFFE", X"FFFD", X"FFFD", X"FFFD", X"FFFD", 
X"FFFD", X"FFFD", X"FFFD", X"FFFD", X"FFFC", X"FFFC", X"FFFC", X"FFFC", X"FFFC", X"FFFC", 
X"FFFC", X"FFFB", X"FFFB", X"FFFB", X"FFFB", X"FFFB", X"FFFB", X"FFFB", X"FFFA", X"FFFA", 
X"FFFA", X"FFFA", X"FFFA", X"FFFA", X"FFF9", X"FFF9", X"FFF9", X"FFF9", X"FFF9", X"FFF8", 
X"FFF8", X"FFF8", X"FFF8", X"FFF8", X"FFF7", X"FFF7", X"FFF7", X"FFF7", X"FFF7", X"FFF6", 
X"FFF6", X"FFF6", X"FFF6", X"FFF5", X"FFF5", X"FFF5", X"FFF5", X"FFF5", X"FFF4", X"FFF4", 
X"FFF4", X"FFF4", X"FFF3", X"FFF3", X"FFF3", X"FFF3", X"FFF2", X"FFF2", X"FFF2", X"FFF2", 
X"FFF1", X"FFF1", X"FFF1", X"FFF0", X"FFF0", X"FFF0", X"FFF0", X"FFEF", X"FFEF", X"FFEF", 
X"FFEE", X"FFEE", X"FFEE", X"FFEE", X"FFED", X"FFED", X"FFED", X"FFEC", X"FFEC", X"FFEC", 
X"FFEB", X"FFEB", X"FFEB", X"FFEA", X"FFEA", X"FFEA", X"FFE9", X"FFE9", X"FFE9", X"FFE8", 
X"FFE8", X"FFE8", X"FFE7", X"FFE7", X"FFE7", X"FFE6", X"FFE6", X"FFE6", X"FFE5", X"FFE5", 
X"FFE5", X"FFE4", X"FFE4", X"FFE3", X"FFE3", X"FFE3", X"FFE2", X"FFE2", X"FFE2", X"FFE1", 
X"FFE1", X"FFE0", X"FFE0", X"FFE0", X"FFDF", X"FFDF", X"FFDE", X"FFDE", X"FFDE", X"FFDD", 
X"FFDD", X"FFDC", X"FFDC", X"FFDC", X"FFDB", X"FFDB", X"FFDA", X"FFDA", X"FFD9", X"FFD9", 
X"FFD9", X"FFD8", X"FFD8", X"FFD7", X"FFD7", X"FFD6", X"FFD6", X"FFD5", X"FFD5", X"FFD4", 
X"FFD4", X"FFD4", X"FFD3", X"FFD3", X"FFD2", X"FFD2", X"FFD1", X"FFD1", X"FFD0", X"FFD0", 
X"FFCF", X"FFCF", X"FFCE", X"FFCE", X"FFCD", X"FFCD", X"FFCC", X"FFCC", X"FFCB", X"FFCB", 
X"FFCA", X"FFCA", X"FFC9", X"FFC9", X"FFC8", X"FFC8", X"FFC7", X"FFC7", X"FFC6", X"FFC6", 
X"FFC5", X"FFC5", X"FFC4", X"FFC3", X"FFC3", X"FFC2", X"FFC2", X"FFC1", X"FFC1", X"FFC0", 
X"FFC0", X"FFBF", X"FFBE", X"FFBE", X"FFBD", X"FFBD", X"FFBC", X"FFBC", X"FFBB", X"FFBA", 
X"FFBA", X"FFB9", X"FFB9", X"FFB8", X"FFB7", X"FFB7", X"FFB6", X"FFB6", X"FFB5", X"FFB4", 
X"FFB4", X"FFB3", X"FFB3", X"FFB2", X"FFB1", X"FFB1", X"FFB0", X"FFB0", X"FFAF", X"FFAE", 
X"FFAE", X"FFAD", X"FFAC", X"FFAC", X"FFAB", X"FFAA", X"FFAA", X"FFA9", X"FFA9", X"FFA8", 
X"FFA7", X"FFA7", X"FFA6", X"FFA5", X"FFA5", X"FFA4", X"FFA3", X"FFA3", X"FFA2", X"FFA1", 
X"FFA1", X"FFA0", X"FF9F", X"FF9E", X"FF9E", X"FF9D", X"FF9C", X"FF9C", X"FF9B", X"FF9A", 
X"FF9A", X"FF99", X"FF98", X"FF97", X"FF97", X"FF96", X"FF95", X"FF95", X"FF94", X"FF93", 
X"FF92", X"FF92", X"FF91", X"FF90", X"FF8F", X"FF8F", X"FF8E", X"FF8D", X"FF8C", X"FF8C", 
X"FF8B", X"FF8A", X"FF89", X"FF89", X"FF88", X"FF87", X"FF86", X"FF86", X"FF85", X"FF84", 
X"FF83", X"FF83", X"FF82", X"FF81", X"FF80", X"FF7F", X"FF7F", X"FF7E", X"FF7D", X"FF7C", 
X"FF7B", X"FF7B", X"FF7A", X"FF79", X"FF78", X"FF77", X"FF77", X"FF76", X"FF75", X"FF74", 
X"FF73", X"FF72", X"FF72", X"FF71", X"FF70", X"FF6F", X"FF6E", X"FF6D", X"FF6D", X"FF6C", 
X"FF6B", X"FF6A", X"FF69", X"FF68", X"FF67", X"FF67", X"FF66", X"FF65", X"FF64", X"FF63", 
X"FF62", X"FF61", X"FF60", X"FF60", X"FF5F", X"FF5E", X"FF5D", X"FF5C", X"FF5B", X"FF5A", 
X"FF59", X"FF58", X"FF58", X"FF57", X"FF56", X"FF55", X"FF54", X"FF53", X"FF52", X"FF51", 
X"FF50", X"FF4F", X"FF4E", X"FF4D", X"FF4C", X"FF4C", X"FF4B", X"FF4A", X"FF49", X"FF48", 
X"FF47", X"FF46", X"FF45", X"FF44", X"FF43", X"FF42", X"FF41", X"FF40", X"FF3F", X"FF3E", 
X"FF3D", X"FF3C", X"FF3B", X"FF3A", X"FF39", X"FF38", X"FF37", X"FF36", X"FF35", X"FF34", 
X"FF33", X"FF32", X"FF31", X"FF30", X"FF2F", X"FF2E", X"FF2D", X"FF2C", X"FF2B", X"FF2A", 
X"FF29", X"FF28", X"FF27", X"FF26", X"FF25", X"FF24", X"FF23", X"FF22", X"FF21", X"FF20", 
X"FF1F", X"FF1E", X"FF1D", X"FF1C", X"FF1B", X"FF1A", X"FF19", X"FF18", X"FF17", X"FF15", 
X"FF14", X"FF13", X"FF12", X"FF11", X"FF10", X"FF0F", X"FF0E", X"FF0D", X"FF0C", X"FF0B", 
X"FF0A", X"FF08", X"FF07", X"FF06", X"FF05", X"FF04", X"FF03", X"FF02", X"FF01", X"FF00", 
X"FEFF", X"FEFD", X"FEFC", X"FEFB", X"FEFA", X"FEF9", X"FEF8", X"FEF7", X"FEF5", X"FEF4", 
X"FEF3", X"FEF2", X"FEF1", X"FEF0", X"FEEF", X"FEED", X"FEEC", X"FEEB", X"FEEA", X"FEE9", 
X"FEE8", X"FEE6", X"FEE5", X"FEE4", X"FEE3", X"FEE2", X"FEE1", X"FEDF", X"FEDE", X"FEDD", 
X"FEDC", X"FEDB", X"FED9", X"FED8", X"FED7", X"FED6", X"FED5", X"FED3", X"FED2", X"FED1", 
X"FED0", X"FECF", X"FECD", X"FECC", X"FECB", X"FECA", X"FEC9", X"FEC7", X"FEC6", X"FEC5", 
X"FEC4", X"FEC2", X"FEC1", X"FEC0", X"FEBF", X"FEBD", X"FEBC", X"FEBB", X"FEBA", X"FEB8", 
X"FEB7", X"FEB6", X"FEB5", X"FEB3", X"FEB2", X"FEB1", X"FEAF", X"FEAE", X"FEAD", X"FEAC", 
X"FEAA", X"FEA9", X"FEA8", X"FEA6", X"FEA5", X"FEA4", X"FEA3", X"FEA1", X"FEA0", X"FE9F", 
X"FE9D", X"FE9C", X"FE9B", X"FE99", X"FE98", X"FE97", X"FE95", X"FE94", X"FE93", X"FE91", 
X"FE90", X"FE8F", X"FE8D", X"FE8C", X"FE8B", X"FE89", X"FE88", X"FE87", X"FE85", X"FE84", 
X"FE83", X"FE81", X"FE80", X"FE7F", X"FE7D", X"FE7C", X"FE7A", X"FE79", X"FE78", X"FE76", 
X"FE75", X"FE74", X"FE72", X"FE71", X"FE6F", X"FE6E", X"FE6D", X"FE6B", X"FE6A", X"FE68", 
X"FE67", X"FE66", X"FE64", X"FE63", X"FE61", X"FE60", X"FE5E", X"FE5D", X"FE5C", X"FE5A", 
X"FE59", X"FE57", X"FE56", X"FE54", X"FE53", X"FE52", X"FE50", X"FE4F", X"FE4D", X"FE4C", 
X"FE4A", X"FE49", X"FE47", X"FE46", X"FE44", X"FE43", X"FE42", X"FE40", X"FE3F", X"FE3D", 
X"FE3C", X"FE3A", X"FE39", X"FE37", X"FE36", X"FE34", X"FE33", X"FE31", X"FE30", X"FE2E", 
X"FE2D", X"FE2B", X"FE2A", X"FE28", X"FE27", X"FE25", X"FE24", X"FE22", X"FE21", X"FE1F", 
X"FE1E", X"FE1C", X"FE1B", X"FE19", X"FE17", X"FE16", X"FE14", X"FE13", X"FE11", X"FE10", 
X"FE0E", X"FE0D", X"FE0B", X"FE0A", X"FE08", X"FE06", X"FE05", X"FE03", X"FE02", X"FE00", 
X"FDFF", X"FDFD", X"FDFB", X"FDFA", X"FDF8", X"FDF7", X"FDF5", X"FDF3", X"FDF2", X"FDF0", 
X"FDEF", X"FDED", X"FDEB", X"FDEA", X"FDE8", X"FDE7", X"FDE5", X"FDE3", X"FDE2", X"FDE0", 
X"FDDF", X"FDDD", X"FDDB", X"FDDA", X"FDD8", X"FDD6", X"FDD5", X"FDD3", X"FDD1", X"FDD0", 
X"FDCE", X"FDCD", X"FDCB", X"FDC9", X"FDC8", X"FDC6", X"FDC4", X"FDC3", X"FDC1", X"FDBF", 
X"FDBE", X"FDBC", X"FDBA", X"FDB9", X"FDB7", X"FDB5", X"FDB4", X"FDB2", X"FDB0", X"FDAE", 
X"FDAD", X"FDAB", X"FDA9", X"FDA8", X"FDA6", X"FDA4", X"FDA3", X"FDA1", X"FD9F", X"FD9D", 
X"FD9C", X"FD9A", X"FD98", X"FD97", X"FD95", X"FD93", X"FD91", X"FD90", X"FD8E", X"FD8C", 
X"FD8A", X"FD89", X"FD87", X"FD85", X"FD83", X"FD82", X"FD80", X"FD7E", X"FD7C", X"FD7B", 
X"FD79", X"FD77", X"FD75", X"FD74", X"FD72", X"FD70", X"FD6E", X"FD6C", X"FD6B", X"FD69", 
X"FD67", X"FD65", X"FD63", X"FD62", X"FD60", X"FD5E", X"FD5C", X"FD5A", X"FD59", X"FD57", 
X"FD55", X"FD53", X"FD51", X"FD50", X"FD4E", X"FD4C", X"FD4A", X"FD48", X"FD46", X"FD45", 
X"FD43", X"FD41", X"FD3F", X"FD3D", X"FD3B", X"FD3A", X"FD38", X"FD36", X"FD34", X"FD32", 
X"FD30", X"FD2E", X"FD2C", X"FD2B", X"FD29", X"FD27", X"FD25", X"FD23", X"FD21", X"FD1F", 
X"FD1D", X"FD1C", X"FD1A", X"FD18", X"FD16", X"FD14", X"FD12", X"FD10", X"FD0E", X"FD0C", 
X"FD0A", X"FD09", X"FD07", X"FD05", X"FD03", X"FD01", X"FCFF", X"FCFD", X"FCFB", X"FCF9", 
X"FCF7", X"FCF5", X"FCF3", X"FCF1", X"FCF0", X"FCEE", X"FCEC", X"FCEA", X"FCE8", X"FCE6", 
X"FCE4", X"FCE2", X"FCE0", X"FCDE", X"FCDC", X"FCDA", X"FCD8", X"FCD6", X"FCD4", X"FCD2", 
X"FCD0", X"FCCE", X"FCCC", X"FCCA", X"FCC8", X"FCC6", X"FCC4", X"FCC2", X"FCC0", X"FCBE", 
X"FCBC", X"FCBA", X"FCB8", X"FCB6", X"FCB4", X"FCB2", X"FCB0", X"FCAE", X"FCAC", X"FCAA", 
X"FCA8", X"FCA6", X"FCA4", X"FCA2", X"FCA0", X"FC9E", X"FC9C", X"FC9A", X"FC98", X"FC96", 
X"FC94", X"FC92", X"FC8F", X"FC8D", X"FC8B", X"FC89", X"FC87", X"FC85", X"FC83", X"FC81", 
X"FC7F", X"FC7D", X"FC7B", X"FC79", X"FC77", X"FC75", X"FC72", X"FC70", X"FC6E", X"FC6C", 
X"FC6A", X"FC68", X"FC66", X"FC64", X"FC62", X"FC60", X"FC5D", X"FC5B", X"FC59", X"FC57", 
X"FC55", X"FC53", X"FC51", X"FC4F", X"FC4C", X"FC4A", X"FC48", X"FC46", X"FC44", X"FC42", 
X"FC40", X"FC3D", X"FC3B", X"FC39", X"FC37", X"FC35", X"FC33", X"FC30", X"FC2E", X"FC2C", 
X"FC2A", X"FC28", X"FC26", X"FC23", X"FC21", X"FC1F", X"FC1D", X"FC1B", X"FC19", X"FC16", 
X"FC14", X"FC12", X"FC10", X"FC0E", X"FC0B", X"FC09", X"FC07", X"FC05", X"FC03", X"FC00", 
X"FBFE", X"FBFC", X"FBFA", X"FBF7", X"FBF5", X"FBF3", X"FBF1", X"FBEE", X"FBEC", X"FBEA", 
X"FBE8", X"FBE6", X"FBE3", X"FBE1", X"FBDF", X"FBDD", X"FBDA", X"FBD8", X"FBD6", X"FBD4", 
X"FBD1", X"FBCF", X"FBCD", X"FBCA", X"FBC8", X"FBC6", X"FBC4", X"FBC1", X"FBBF", X"FBBD", 
X"FBBA", X"FBB8", X"FBB6", X"FBB4", X"FBB1", X"FBAF", X"FBAD", X"FBAA", X"FBA8", X"FBA6", 
X"FBA3", X"FBA1", X"FB9F", X"FB9D", X"FB9A", X"FB98", X"FB96", X"FB93", X"FB91", X"FB8F", 
X"FB8C", X"FB8A", X"FB88", X"FB85", X"FB83", X"FB81", X"FB7E", X"FB7C", X"FB79", X"FB77", 
X"FB75", X"FB72", X"FB70", X"FB6E", X"FB6B", X"FB69", X"FB67", X"FB64", X"FB62", X"FB5F", 
X"FB5D", X"FB5B", X"FB58", X"FB56", X"FB53", X"FB51", X"FB4F", X"FB4C", X"FB4A", X"FB47", 
X"FB45", X"FB43", X"FB40", X"FB3E", X"FB3B", X"FB39", X"FB37", X"FB34", X"FB32", X"FB2F", 
X"FB2D", X"FB2A", X"FB28", X"FB26", X"FB23", X"FB21", X"FB1E", X"FB1C", X"FB19", X"FB17", 
X"FB14", X"FB12", X"FB10", X"FB0D", X"FB0B", X"FB08", X"FB06", X"FB03", X"FB01", X"FAFE", 
X"FAFC", X"FAF9", X"FAF7", X"FAF4", X"FAF2", X"FAEF", X"FAED", X"FAEA", X"FAE8", X"FAE5", 
X"FAE3", X"FAE0", X"FADE", X"FADB", X"FAD9", X"FAD6", X"FAD4", X"FAD1", X"FACF", X"FACC", 
X"FACA", X"FAC7", X"FAC5", X"FAC2", X"FAC0", X"FABD", X"FABB", X"FAB8", X"FAB6", X"FAB3", 
X"FAB0", X"FAAE", X"FAAB", X"FAA9", X"FAA6", X"FAA4", X"FAA1", X"FA9F", X"FA9C", X"FA99", 
X"FA97", X"FA94", X"FA92", X"FA8F", X"FA8D", X"FA8A", X"FA87", X"FA85", X"FA82", X"FA80", 
X"FA7D", X"FA7A", X"FA78", X"FA75", X"FA73", X"FA70", X"FA6D", X"FA6B", X"FA68", X"FA66", 
X"FA63", X"FA60", X"FA5E", X"FA5B", X"FA58", X"FA56", X"FA53", X"FA51", X"FA4E", X"FA4B", 
X"FA49", X"FA46", X"FA43", X"FA41", X"FA3E", X"FA3B", X"FA39", X"FA36", X"FA33", X"FA31", 
X"FA2E", X"FA2B", X"FA29", X"FA26", X"FA23", X"FA21", X"FA1E", X"FA1B", X"FA19", X"FA16", 
X"FA13", X"FA11", X"FA0E", X"FA0B", X"FA09", X"FA06", X"FA03", X"FA01", X"F9FE", X"F9FB", 
X"F9F8", X"F9F6", X"F9F3", X"F9F0", X"F9EE", X"F9EB", X"F9E8", X"F9E5", X"F9E3", X"F9E0", 
X"F9DD", X"F9DA", X"F9D8", X"F9D5", X"F9D2", X"F9CF", X"F9CD", X"F9CA", X"F9C7", X"F9C4", 
X"F9C2", X"F9BF", X"F9BC", X"F9B9", X"F9B7", X"F9B4", X"F9B1", X"F9AE", X"F9AC", X"F9A9", 
X"F9A6", X"F9A3", X"F9A0", X"F99E", X"F99B", X"F998", X"F995", X"F993", X"F990", X"F98D", 
X"F98A", X"F987", X"F985", X"F982", X"F97F", X"F97C", X"F979", X"F976", X"F974", X"F971", 
X"F96E", X"F96B", X"F968", X"F966", X"F963", X"F960", X"F95D", X"F95A", X"F957", X"F954", 
X"F952", X"F94F", X"F94C", X"F949", X"F946", X"F943", X"F940", X"F93E", X"F93B", X"F938", 
X"F935", X"F932", X"F92F", X"F92C", X"F929", X"F927", X"F924", X"F921", X"F91E", X"F91B", 
X"F918", X"F915", X"F912", X"F90F", X"F90D", X"F90A", X"F907", X"F904", X"F901", X"F8FE", 
X"F8FB", X"F8F8", X"F8F5", X"F8F2", X"F8EF", X"F8EC", X"F8EA", X"F8E7", X"F8E4", X"F8E1", 
X"F8DE", X"F8DB", X"F8D8", X"F8D5", X"F8D2", X"F8CF", X"F8CC", X"F8C9", X"F8C6", X"F8C3", 
X"F8C0", X"F8BD", X"F8BA", X"F8B7", X"F8B4", X"F8B1", X"F8AE", X"F8AB", X"F8A8", X"F8A5", 
X"F8A3", X"F8A0", X"F89D", X"F89A", X"F897", X"F894", X"F891", X"F88E", X"F88B", X"F888", 
X"F885", X"F882", X"F87E", X"F87B", X"F878", X"F875", X"F872", X"F86F", X"F86C", X"F869", 
X"F866", X"F863", X"F860", X"F85D", X"F85A", X"F857", X"F854", X"F851", X"F84E", X"F84B", 
X"F848", X"F845", X"F842", X"F83F", X"F83C", X"F839", X"F835", X"F832", X"F82F", X"F82C", 
X"F829", X"F826", X"F823", X"F820", X"F81D", X"F81A", X"F817", X"F814", X"F810", X"F80D", 
X"F80A", X"F807", X"F804", X"F801", X"F7FE", X"F7FB", X"F7F8", X"F7F4", X"F7F1", X"F7EE", 
X"F7EB", X"F7E8", X"F7E5", X"F7E2", X"F7DF", X"F7DB", X"F7D8", X"F7D5", X"F7D2", X"F7CF", 
X"F7CC", X"F7C9", X"F7C5", X"F7C2", X"F7BF", X"F7BC", X"F7B9", X"F7B6", X"F7B3", X"F7AF", 
X"F7AC", X"F7A9", X"F7A6", X"F7A3", X"F79F", X"F79C", X"F799", X"F796", X"F793", X"F790", 
X"F78C", X"F789", X"F786", X"F783", X"F780", X"F77C", X"F779", X"F776", X"F773", X"F770", 
X"F76C", X"F769", X"F766", X"F763", X"F75F", X"F75C", X"F759", X"F756", X"F753", X"F74F", 
X"F74C", X"F749", X"F746", X"F742", X"F73F", X"F73C", X"F739", X"F735", X"F732", X"F72F", 
X"F72C", X"F728", X"F725", X"F722", X"F71E", X"F71B", X"F718", X"F715", X"F711", X"F70E", 
X"F70B", X"F708", X"F704", X"F701", X"F6FE", X"F6FA", X"F6F7", X"F6F4", X"F6F0", X"F6ED", 
X"F6EA", X"F6E7", X"F6E3", X"F6E0", X"F6DD", X"F6D9", X"F6D6", X"F6D3", X"F6CF", X"F6CC", 
X"F6C9", X"F6C5", X"F6C2", X"F6BF", X"F6BB", X"F6B8", X"F6B5", X"F6B1", X"F6AE", X"F6AB", 
X"F6A7", X"F6A4", X"F6A1", X"F69D", X"F69A", X"F696", X"F693", X"F690", X"F68C", X"F689", 
X"F686", X"F682", X"F67F", X"F67B", X"F678", X"F675", X"F671", X"F66E", X"F66B", X"F667", 
X"F664", X"F660", X"F65D", X"F65A", X"F656", X"F653", X"F64F", X"F64C", X"F649", X"F645", 
X"F642", X"F63E", X"F63B", X"F637", X"F634", X"F631", X"F62D", X"F62A", X"F626", X"F623", 
X"F61F", X"F61C", X"F618", X"F615", X"F612", X"F60E", X"F60B", X"F607", X"F604", X"F600", 
X"F5FD", X"F5F9", X"F5F6", X"F5F2", X"F5EF", X"F5EB", X"F5E8", X"F5E5", X"F5E1", X"F5DE", 
X"F5DA", X"F5D7", X"F5D3", X"F5D0", X"F5CC", X"F5C9", X"F5C5", X"F5C2", X"F5BE", X"F5BB", 
X"F5B7", X"F5B4", X"F5B0", X"F5AD", X"F5A9", X"F5A6", X"F5A2", X"F59E", X"F59B", X"F597", 
X"F594", X"F590", X"F58D", X"F589", X"F586", X"F582", X"F57F", X"F57B", X"F578", X"F574", 
X"F570", X"F56D", X"F569", X"F566", X"F562", X"F55F", X"F55B", X"F558", X"F554", X"F550", 
X"F54D", X"F549", X"F546", X"F542", X"F53E", X"F53B", X"F537", X"F534", X"F530", X"F52D", 
X"F529", X"F525", X"F522", X"F51E", X"F51B", X"F517", X"F513", X"F510", X"F50C", X"F508", 
X"F505", X"F501", X"F4FE", X"F4FA", X"F4F6", X"F4F3", X"F4EF", X"F4EB", X"F4E8", X"F4E4", 
X"F4E1", X"F4DD", X"F4D9", X"F4D6", X"F4D2", X"F4CE", X"F4CB", X"F4C7", X"F4C3", X"F4C0", 
X"F4BC", X"F4B8", X"F4B5", X"F4B1", X"F4AD", X"F4AA", X"F4A6", X"F4A2", X"F49F", X"F49B", 
X"F497", X"F493", X"F490", X"F48C", X"F488", X"F485", X"F481", X"F47D", X"F47A", X"F476", 
X"F472", X"F46E", X"F46B", X"F467", X"F463", X"F460", X"F45C", X"F458", X"F454", X"F451", 
X"F44D", X"F449", X"F446", X"F442", X"F43E", X"F43A", X"F437", X"F433", X"F42F", X"F42B", 
X"F428", X"F424", X"F420", X"F41C", X"F419", X"F415", X"F411", X"F40D", X"F409", X"F406", 
X"F402", X"F3FE", X"F3FA", X"F3F7", X"F3F3", X"F3EF", X"F3EB", X"F3E7", X"F3E4", X"F3E0", 
X"F3DC", X"F3D8", X"F3D4", X"F3D1", X"F3CD", X"F3C9", X"F3C5", X"F3C1", X"F3BE", X"F3BA", 
X"F3B6", X"F3B2", X"F3AE", X"F3AA", X"F3A7", X"F3A3", X"F39F", X"F39B", X"F397", X"F393", 
X"F390", X"F38C", X"F388", X"F384", X"F380", X"F37C", X"F379", X"F375", X"F371", X"F36D", 
X"F369", X"F365", X"F361", X"F35D", X"F35A", X"F356", X"F352", X"F34E", X"F34A", X"F346", 
X"F342", X"F33E", X"F33B", X"F337", X"F333", X"F32F", X"F32B", X"F327", X"F323", X"F31F", 
X"F31B", X"F317", X"F314", X"F310", X"F30C", X"F308", X"F304", X"F300", X"F2FC", X"F2F8", 
X"F2F4", X"F2F0", X"F2EC", X"F2E8", X"F2E4", X"F2E0", X"F2DD", X"F2D9", X"F2D5", X"F2D1", 
X"F2CD", X"F2C9", X"F2C5", X"F2C1", X"F2BD", X"F2B9", X"F2B5", X"F2B1", X"F2AD", X"F2A9", 
X"F2A5", X"F2A1", X"F29D", X"F299", X"F295", X"F291", X"F28D", X"F289", X"F285", X"F281", 
X"F27D", X"F279", X"F275", X"F271", X"F26D", X"F269", X"F265", X"F261", X"F25D", X"F259", 
X"F255", X"F251", X"F24D", X"F249", X"F245", X"F241", X"F23D", X"F239", X"F235", X"F231", 
X"F22D", X"F229", X"F225", X"F221", X"F21D", X"F219", X"F215", X"F211", X"F20D", X"F208", 
X"F204", X"F200", X"F1FC", X"F1F8", X"F1F4", X"F1F0", X"F1EC", X"F1E8", X"F1E4", X"F1E0", 
X"F1DC", X"F1D8", X"F1D3", X"F1CF", X"F1CB", X"F1C7", X"F1C3", X"F1BF", X"F1BB", X"F1B7", 
X"F1B3", X"F1AF", X"F1AB", X"F1A6", X"F1A2", X"F19E", X"F19A", X"F196", X"F192", X"F18E", 
X"F18A", X"F185", X"F181", X"F17D", X"F179", X"F175", X"F171", X"F16D", X"F168", X"F164", 
X"F160", X"F15C", X"F158", X"F154", X"F150", X"F14B", X"F147", X"F143", X"F13F", X"F13B", 
X"F137", X"F132", X"F12E", X"F12A", X"F126", X"F122", X"F11E", X"F119", X"F115", X"F111", 
X"F10D", X"F109", X"F104", X"F100", X"F0FC", X"F0F8", X"F0F4", X"F0EF", X"F0EB", X"F0E7", 
X"F0E3", X"F0DF", X"F0DA", X"F0D6", X"F0D2", X"F0CE", X"F0C9", X"F0C5", X"F0C1", X"F0BD", 
X"F0B9", X"F0B4", X"F0B0", X"F0AC", X"F0A8", X"F0A3", X"F09F", X"F09B", X"F097", X"F092", 
X"F08E", X"F08A", X"F086", X"F081", X"F07D", X"F079", X"F075", X"F070", X"F06C", X"F068", 
X"F063", X"F05F", X"F05B", X"F057", X"F052", X"F04E", X"F04A", X"F045", X"F041", X"F03D", 
X"F039", X"F034", X"F030", X"F02C", X"F027", X"F023", X"F01F", X"F01A", X"F016", X"F012", 
X"F00D", X"F009", X"F005", X"F001", X"EFFC", X"EFF8", X"EFF4", X"EFEF", X"EFEB", X"EFE7", 
X"EFE2", X"EFDE", X"EFDA", X"EFD5", X"EFD1", X"EFCC", X"EFC8", X"EFC4", X"EFBF", X"EFBB", 
X"EFB7", X"EFB2", X"EFAE", X"EFAA", X"EFA5", X"EFA1", X"EF9C", X"EF98", X"EF94", X"EF8F", 
X"EF8B", X"EF87", X"EF82", X"EF7E", X"EF79", X"EF75", X"EF71", X"EF6C", X"EF68", X"EF63", 
X"EF5F", X"EF5B", X"EF56", X"EF52", X"EF4D", X"EF49", X"EF45", X"EF40", X"EF3C", X"EF37", 
X"EF33", X"EF2E", X"EF2A", X"EF26", X"EF21", X"EF1D", X"EF18", X"EF14", X"EF0F", X"EF0B", 
X"EF06", X"EF02", X"EEFE", X"EEF9", X"EEF5", X"EEF0", X"EEEC", X"EEE7", X"EEE3", X"EEDE", 
X"EEDA", X"EED5", X"EED1", X"EECD", X"EEC8", X"EEC4", X"EEBF", X"EEBB", X"EEB6", X"EEB2", 
X"EEAD", X"EEA9", X"EEA4", X"EEA0", X"EE9B", X"EE97", X"EE92", X"EE8E", X"EE89", X"EE85", 
X"EE80", X"EE7C", X"EE77", X"EE73", X"EE6E", X"EE6A", X"EE65", X"EE61", X"EE5C", X"EE57", 
X"EE53", X"EE4E", X"EE4A", X"EE45", X"EE41", X"EE3C", X"EE38", X"EE33", X"EE2F", X"EE2A", 
X"EE26", X"EE21", X"EE1C", X"EE18", X"EE13", X"EE0F", X"EE0A", X"EE06", X"EE01", X"EDFC", 
X"EDF8", X"EDF3", X"EDEF", X"EDEA", X"EDE6", X"EDE1", X"EDDC", X"EDD8", X"EDD3", X"EDCF", 
X"EDCA", X"EDC5", X"EDC1", X"EDBC", X"EDB8", X"EDB3", X"EDAE", X"EDAA", X"EDA5", X"EDA1", 
X"ED9C", X"ED97", X"ED93", X"ED8E", X"ED8A", X"ED85", X"ED80", X"ED7C", X"ED77", X"ED72", 
X"ED6E", X"ED69", X"ED64", X"ED60", X"ED5B", X"ED57", X"ED52", X"ED4D", X"ED49", X"ED44", 
X"ED3F", X"ED3B", X"ED36", X"ED31", X"ED2D", X"ED28", X"ED23", X"ED1F", X"ED1A", X"ED15", 
X"ED11", X"ED0C", X"ED07", X"ED03", X"ECFE", X"ECF9", X"ECF5", X"ECF0", X"ECEB", X"ECE6", 
X"ECE2", X"ECDD", X"ECD8", X"ECD4", X"ECCF", X"ECCA", X"ECC6", X"ECC1", X"ECBC", X"ECB7", 
X"ECB3", X"ECAE", X"ECA9", X"ECA4", X"ECA0", X"EC9B", X"EC96", X"EC92", X"EC8D", X"EC88", 
X"EC83", X"EC7F", X"EC7A", X"EC75", X"EC70", X"EC6C", X"EC67", X"EC62", X"EC5D", X"EC59", 
X"EC54", X"EC4F", X"EC4A", X"EC46", X"EC41", X"EC3C", X"EC37", X"EC32", X"EC2E", X"EC29", 
X"EC24", X"EC1F", X"EC1B", X"EC16", X"EC11", X"EC0C", X"EC07", X"EC03", X"EBFE", X"EBF9", 
X"EBF4", X"EBEF", X"EBEB", X"EBE6", X"EBE1", X"EBDC", X"EBD7", X"EBD3", X"EBCE", X"EBC9", 
X"EBC4", X"EBBF", X"EBBA", X"EBB6", X"EBB1", X"EBAC", X"EBA7", X"EBA2", X"EB9D", X"EB99", 
X"EB94", X"EB8F", X"EB8A", X"EB85", X"EB80", X"EB7C", X"EB77", X"EB72", X"EB6D", X"EB68", 
X"EB63", X"EB5E", X"EB5A", X"EB55", X"EB50", X"EB4B", X"EB46", X"EB41", X"EB3C", X"EB37", 
X"EB33", X"EB2E", X"EB29", X"EB24", X"EB1F", X"EB1A", X"EB15", X"EB10", X"EB0B", X"EB07", 
X"EB02", X"EAFD", X"EAF8", X"EAF3", X"EAEE", X"EAE9", X"EAE4", X"EADF", X"EADA", X"EAD5", 
X"EAD0", X"EACC", X"EAC7", X"EAC2", X"EABD", X"EAB8", X"EAB3", X"EAAE", X"EAA9", X"EAA4", 
X"EA9F", X"EA9A", X"EA95", X"EA90", X"EA8B", X"EA86", X"EA81", X"EA7C", X"EA78", X"EA73", 
X"EA6E", X"EA69", X"EA64", X"EA5F", X"EA5A", X"EA55", X"EA50", X"EA4B", X"EA46", X"EA41", 
X"EA3C", X"EA37", X"EA32", X"EA2D", X"EA28", X"EA23", X"EA1E", X"EA19", X"EA14", X"EA0F", 
X"EA0A", X"EA05", X"EA00", X"E9FB", X"E9F6", X"E9F1", X"E9EC", X"E9E7", X"E9E2", X"E9DD", 
X"E9D8", X"E9D3", X"E9CE", X"E9C9", X"E9C4", X"E9BF", X"E9BA", X"E9B5", X"E9AF", X"E9AA", 
X"E9A5", X"E9A0", X"E99B", X"E996", X"E991", X"E98C", X"E987", X"E982", X"E97D", X"E978", 
X"E973", X"E96E", X"E969", X"E964", X"E95F", X"E959", X"E954", X"E94F", X"E94A", X"E945", 
X"E940", X"E93B", X"E936", X"E931", X"E92C", X"E927", X"E922", X"E91C", X"E917", X"E912", 
X"E90D", X"E908", X"E903", X"E8FE", X"E8F9", X"E8F4", X"E8EE", X"E8E9", X"E8E4", X"E8DF", 
X"E8DA", X"E8D5", X"E8D0", X"E8CB", X"E8C5", X"E8C0", X"E8BB", X"E8B6", X"E8B1", X"E8AC", 
X"E8A7", X"E8A1", X"E89C", X"E897", X"E892", X"E88D", X"E888", X"E883", X"E87D", X"E878", 
X"E873", X"E86E", X"E869", X"E864", X"E85E", X"E859", X"E854", X"E84F", X"E84A", X"E844", 
X"E83F", X"E83A", X"E835", X"E830", X"E82B", X"E825", X"E820", X"E81B", X"E816", X"E811", 
X"E80B", X"E806", X"E801", X"E7FC", X"E7F7", X"E7F1", X"E7EC", X"E7E7", X"E7E2", X"E7DC", 
X"E7D7", X"E7D2", X"E7CD", X"E7C8", X"E7C2", X"E7BD", X"E7B8", X"E7B3", X"E7AD", X"E7A8", 
X"E7A3", X"E79E", X"E798", X"E793", X"E78E", X"E789", X"E783", X"E77E", X"E779", X"E774", 
X"E76E", X"E769", X"E764", X"E75F", X"E759", X"E754", X"E74F", X"E749", X"E744", X"E73F", 
X"E73A", X"E734", X"E72F", X"E72A", X"E724", X"E71F", X"E71A", X"E715", X"E70F", X"E70A", 
X"E705", X"E6FF", X"E6FA", X"E6F5", X"E6EF", X"E6EA", X"E6E5", X"E6DF", X"E6DA", X"E6D5", 
X"E6D0", X"E6CA", X"E6C5", X"E6C0", X"E6BA", X"E6B5", X"E6B0", X"E6AA", X"E6A5", X"E6A0", 
X"E69A", X"E695", X"E68F", X"E68A", X"E685", X"E67F", X"E67A", X"E675", X"E66F", X"E66A", 
X"E665", X"E65F", X"E65A", X"E655", X"E64F", X"E64A", X"E644", X"E63F", X"E63A", X"E634", 
X"E62F", X"E62A", X"E624", X"E61F", X"E619", X"E614", X"E60F", X"E609", X"E604", X"E5FE", 
X"E5F9", X"E5F4", X"E5EE", X"E5E9", X"E5E3", X"E5DE", X"E5D9", X"E5D3", X"E5CE", X"E5C8", 
X"E5C3", X"E5BD", X"E5B8", X"E5B3", X"E5AD", X"E5A8", X"E5A2", X"E59D", X"E597", X"E592", 
X"E58D", X"E587", X"E582", X"E57C", X"E577", X"E571", X"E56C", X"E566", X"E561", X"E55C", 
X"E556", X"E551", X"E54B", X"E546", X"E540", X"E53B", X"E535", X"E530", X"E52A", X"E525", 
X"E51F", X"E51A", X"E514", X"E50F", X"E509", X"E504", X"E4FF", X"E4F9", X"E4F4", X"E4EE", 
X"E4E9", X"E4E3", X"E4DE", X"E4D8", X"E4D3", X"E4CD", X"E4C8", X"E4C2", X"E4BC", X"E4B7", 
X"E4B1", X"E4AC", X"E4A6", X"E4A1", X"E49B", X"E496", X"E490", X"E48B", X"E485", X"E480", 
X"E47A", X"E475", X"E46F", X"E46A", X"E464", X"E45E", X"E459", X"E453", X"E44E", X"E448", 
X"E443", X"E43D", X"E438", X"E432", X"E42D", X"E427", X"E421", X"E41C", X"E416", X"E411", 
X"E40B", X"E406", X"E400", X"E3FA", X"E3F5", X"E3EF", X"E3EA", X"E3E4", X"E3DE", X"E3D9", 
X"E3D3", X"E3CE", X"E3C8", X"E3C2", X"E3BD", X"E3B7", X"E3B2", X"E3AC", X"E3A6", X"E3A1", 
X"E39B", X"E396", X"E390", X"E38A", X"E385", X"E37F", X"E37A", X"E374", X"E36E", X"E369", 
X"E363", X"E35D", X"E358", X"E352", X"E34C", X"E347", X"E341", X"E33C", X"E336", X"E330", 
X"E32B", X"E325", X"E31F", X"E31A", X"E314", X"E30E", X"E309", X"E303", X"E2FD", X"E2F8", 
X"E2F2", X"E2EC", X"E2E7", X"E2E1", X"E2DB", X"E2D6", X"E2D0", X"E2CA", X"E2C5", X"E2BF", 
X"E2B9", X"E2B4", X"E2AE", X"E2A8", X"E2A2", X"E29D", X"E297", X"E291", X"E28C", X"E286", 
X"E280", X"E27B", X"E275", X"E26F", X"E269", X"E264", X"E25E", X"E258", X"E253", X"E24D", 
X"E247", X"E241", X"E23C", X"E236", X"E230", X"E22A", X"E225", X"E21F", X"E219", X"E213", 
X"E20E", X"E208", X"E202", X"E1FD", X"E1F7", X"E1F1", X"E1EB", X"E1E5", X"E1E0", X"E1DA", 
X"E1D4", X"E1CE", X"E1C9", X"E1C3", X"E1BD", X"E1B7", X"E1B2", X"E1AC", X"E1A6", X"E1A0", 
X"E19A", X"E195", X"E18F", X"E189", X"E183", X"E17E", X"E178", X"E172", X"E16C", X"E166", 
X"E161", X"E15B", X"E155", X"E14F", X"E149", X"E144", X"E13E", X"E138", X"E132", X"E12C", 
X"E126", X"E121", X"E11B", X"E115", X"E10F", X"E109", X"E104", X"E0FE", X"E0F8", X"E0F2", 
X"E0EC", X"E0E6", X"E0E1", X"E0DB", X"E0D5", X"E0CF", X"E0C9", X"E0C3", X"E0BD", X"E0B8", 
X"E0B2", X"E0AC", X"E0A6", X"E0A0", X"E09A", X"E094", X"E08F", X"E089", X"E083", X"E07D", 
X"E077", X"E071", X"E06B", X"E065", X"E060", X"E05A", X"E054", X"E04E", X"E048", X"E042", 
X"E03C", X"E036", X"E031", X"E02B", X"E025", X"E01F", X"E019", X"E013", X"E00D", X"E007", 
X"E001", X"DFFB", X"DFF5", X"DFF0", X"DFEA", X"DFE4", X"DFDE", X"DFD8", X"DFD2", X"DFCC", 
X"DFC6", X"DFC0", X"DFBA", X"DFB4", X"DFAE", X"DFA8", X"DFA2", X"DF9D", X"DF97", X"DF91", 
X"DF8B", X"DF85", X"DF7F", X"DF79", X"DF73", X"DF6D", X"DF67", X"DF61", X"DF5B", X"DF55", 
X"DF4F", X"DF49", X"DF43", X"DF3D", X"DF37", X"DF31", X"DF2B", X"DF25", X"DF1F", X"DF19", 
X"DF13", X"DF0D", X"DF07", X"DF01", X"DEFB", X"DEF5", X"DEEF", X"DEE9", X"DEE3", X"DEDD", 
X"DED7", X"DED1", X"DECB", X"DEC5", X"DEBF", X"DEB9", X"DEB3", X"DEAD", X"DEA7", X"DEA1", 
X"DE9B", X"DE95", X"DE8F", X"DE89", X"DE83", X"DE7D", X"DE77", X"DE71", X"DE6B", X"DE65", 
X"DE5F", X"DE59", X"DE53", X"DE4D", X"DE47", X"DE41", X"DE3B", X"DE35", X"DE2F", X"DE29", 
X"DE23", X"DE1D", X"DE17", X"DE10", X"DE0A", X"DE04", X"DDFE", X"DDF8", X"DDF2", X"DDEC", 
X"DDE6", X"DDE0", X"DDDA", X"DDD4", X"DDCE", X"DDC8", X"DDC2", X"DDBB", X"DDB5", X"DDAF", 
X"DDA9", X"DDA3", X"DD9D", X"DD97", X"DD91", X"DD8B", X"DD85", X"DD7F", X"DD78", X"DD72", 
X"DD6C", X"DD66", X"DD60", X"DD5A", X"DD54", X"DD4E", X"DD48", X"DD41", X"DD3B", X"DD35", 
X"DD2F", X"DD29", X"DD23", X"DD1D", X"DD16", X"DD10", X"DD0A", X"DD04", X"DCFE", X"DCF8", 
X"DCF2", X"DCEC", X"DCE5", X"DCDF", X"DCD9", X"DCD3", X"DCCD", X"DCC7", X"DCC0", X"DCBA", 
X"DCB4", X"DCAE", X"DCA8", X"DCA2", X"DC9B", X"DC95", X"DC8F", X"DC89", X"DC83", X"DC7D", 
X"DC76", X"DC70", X"DC6A", X"DC64", X"DC5E", X"DC58", X"DC51", X"DC4B", X"DC45", X"DC3F", 
X"DC39", X"DC32", X"DC2C", X"DC26", X"DC20", X"DC1A", X"DC13", X"DC0D", X"DC07", X"DC01", 
X"DBFA", X"DBF4", X"DBEE", X"DBE8", X"DBE2", X"DBDB", X"DBD5", X"DBCF", X"DBC9", X"DBC2", 
X"DBBC", X"DBB6", X"DBB0", X"DBAA", X"DBA3", X"DB9D", X"DB97", X"DB91", X"DB8A", X"DB84", 
X"DB7E", X"DB78", X"DB71", X"DB6B", X"DB65", X"DB5F", X"DB58", X"DB52", X"DB4C", X"DB46", 
X"DB3F", X"DB39", X"DB33", X"DB2C", X"DB26", X"DB20", X"DB1A", X"DB13", X"DB0D", X"DB07", 
X"DB01", X"DAFA", X"DAF4", X"DAEE", X"DAE7", X"DAE1", X"DADB", X"DAD4", X"DACE", X"DAC8", 
X"DAC2", X"DABB", X"DAB5", X"DAAF", X"DAA8", X"DAA2", X"DA9C", X"DA95", X"DA8F", X"DA89", 
X"DA82", X"DA7C", X"DA76", X"DA70", X"DA69", X"DA63", X"DA5D", X"DA56", X"DA50", X"DA4A", 
X"DA43", X"DA3D", X"DA37", X"DA30", X"DA2A", X"DA24", X"DA1D", X"DA17", X"DA10", X"DA0A", 
X"DA04", X"D9FD", X"D9F7", X"D9F1", X"D9EA", X"D9E4", X"D9DE", X"D9D7", X"D9D1", X"D9CB", 
X"D9C4", X"D9BE", X"D9B7", X"D9B1", X"D9AB", X"D9A4", X"D99E", X"D998", X"D991", X"D98B", 
X"D984", X"D97E", X"D978", X"D971", X"D96B", X"D964", X"D95E", X"D958", X"D951", X"D94B", 
X"D944", X"D93E", X"D938", X"D931", X"D92B", X"D924", X"D91E", X"D918", X"D911", X"D90B", 
X"D904", X"D8FE", X"D8F7", X"D8F1", X"D8EB", X"D8E4", X"D8DE", X"D8D7", X"D8D1", X"D8CA", 
X"D8C4", X"D8BE", X"D8B7", X"D8B1", X"D8AA", X"D8A4", X"D89D", X"D897", X"D890", X"D88A", 
X"D884", X"D87D", X"D877", X"D870", X"D86A", X"D863", X"D85D", X"D856", X"D850", X"D849", 
X"D843", X"D83C", X"D836", X"D82F", X"D829", X"D822", X"D81C", X"D816", X"D80F", X"D809", 
X"D802", X"D7FC", X"D7F5", X"D7EF", X"D7E8", X"D7E2", X"D7DB", X"D7D5", X"D7CE", X"D7C8", 
X"D7C1", X"D7BB", X"D7B4", X"D7AE", X"D7A7", X"D7A1", X"D79A", X"D794", X"D78D", X"D786", 
X"D780", X"D779", X"D773", X"D76C", X"D766", X"D75F", X"D759", X"D752", X"D74C", X"D745", 
X"D73F", X"D738", X"D732", X"D72B", X"D724", X"D71E", X"D717", X"D711", X"D70A", X"D704", 
X"D6FD", X"D6F7", X"D6F0", X"D6EA", X"D6E3", X"D6DC", X"D6D6", X"D6CF", X"D6C9", X"D6C2", 
X"D6BC", X"D6B5", X"D6AE", X"D6A8", X"D6A1", X"D69B", X"D694", X"D68D", X"D687", X"D680", 
X"D67A", X"D673", X"D66D", X"D666", X"D65F", X"D659", X"D652", X"D64C", X"D645", X"D63E", 
X"D638", X"D631", X"D62B", X"D624", X"D61D", X"D617", X"D610", X"D60A", X"D603", X"D5FC", 
X"D5F6", X"D5EF", X"D5E8", X"D5E2", X"D5DB", X"D5D5", X"D5CE", X"D5C7", X"D5C1", X"D5BA", 
X"D5B3", X"D5AD", X"D5A6", X"D59F", X"D599", X"D592", X"D58B", X"D585", X"D57E", X"D578", 
X"D571", X"D56A", X"D564", X"D55D", X"D556", X"D550", X"D549", X"D542", X"D53C", X"D535", 
X"D52E", X"D528", X"D521", X"D51A", X"D514", X"D50D", X"D506", X"D500", X"D4F9", X"D4F2", 
X"D4EB", X"D4E5", X"D4DE", X"D4D7", X"D4D1", X"D4CA", X"D4C3", X"D4BD", X"D4B6", X"D4AF", 
X"D4A9", X"D4A2", X"D49B", X"D494", X"D48E", X"D487", X"D480", X"D47A", X"D473", X"D46C", 
X"D465", X"D45F", X"D458", X"D451", X"D44B", X"D444", X"D43D", X"D436", X"D430", X"D429", 
X"D422", X"D41B", X"D415", X"D40E", X"D407", X"D400", X"D3FA", X"D3F3", X"D3EC", X"D3E6", 
X"D3DF", X"D3D8", X"D3D1", X"D3CA", X"D3C4", X"D3BD", X"D3B6", X"D3AF", X"D3A9", X"D3A2", 
X"D39B", X"D394", X"D38E", X"D387", X"D380", X"D379", X"D373", X"D36C", X"D365", X"D35E", 
X"D357", X"D351", X"D34A", X"D343", X"D33C", X"D335", X"D32F", X"D328", X"D321", X"D31A", 
X"D314", X"D30D", X"D306", X"D2FF", X"D2F8", X"D2F2", X"D2EB", X"D2E4", X"D2DD", X"D2D6", 
X"D2CF", X"D2C9", X"D2C2", X"D2BB", X"D2B4", X"D2AD", X"D2A7", X"D2A0", X"D299", X"D292", 
X"D28B", X"D284", X"D27E", X"D277", X"D270", X"D269", X"D262", X"D25B", X"D255", X"D24E", 
X"D247", X"D240", X"D239", X"D232", X"D22B", X"D225", X"D21E", X"D217", X"D210", X"D209", 
X"D202", X"D1FB", X"D1F5", X"D1EE", X"D1E7", X"D1E0", X"D1D9", X"D1D2", X"D1CB", X"D1C5", 
X"D1BE", X"D1B7", X"D1B0", X"D1A9", X"D1A2", X"D19B", X"D194", X"D18D", X"D187", X"D180", 
X"D179", X"D172", X"D16B", X"D164", X"D15D", X"D156", X"D14F", X"D149", X"D142", X"D13B", 
X"D134", X"D12D", X"D126", X"D11F", X"D118", X"D111", X"D10A", X"D103", X"D0FC", X"D0F6", 
X"D0EF", X"D0E8", X"D0E1", X"D0DA", X"D0D3", X"D0CC", X"D0C5", X"D0BE", X"D0B7", X"D0B0", 
X"D0A9", X"D0A2", X"D09B", X"D095", X"D08E", X"D087", X"D080", X"D079", X"D072", X"D06B", 
X"D064", X"D05D", X"D056", X"D04F", X"D048", X"D041", X"D03A", X"D033", X"D02C", X"D025", 
X"D01E", X"D017", X"D010", X"D009", X"D002", X"CFFB", X"CFF4", X"CFED", X"CFE6", X"CFDF", 
X"CFD8", X"CFD2", X"CFCB", X"CFC4", X"CFBD", X"CFB6", X"CFAF", X"CFA8", X"CFA1", X"CF9A", 
X"CF93", X"CF8C", X"CF85", X"CF7E", X"CF77", X"CF70", X"CF69", X"CF62", X"CF5B", X"CF54", 
X"CF4D", X"CF45", X"CF3E", X"CF37", X"CF30", X"CF29", X"CF22", X"CF1B", X"CF14", X"CF0D", 
X"CF06", X"CEFF", X"CEF8", X"CEF1", X"CEEA", X"CEE3", X"CEDC", X"CED5", X"CECE", X"CEC7", 
X"CEC0", X"CEB9", X"CEB2", X"CEAB", X"CEA4", X"CE9D", X"CE96", X"CE8F", X"CE88", X"CE80", 
X"CE79", X"CE72", X"CE6B", X"CE64", X"CE5D", X"CE56", X"CE4F", X"CE48", X"CE41", X"CE3A", 
X"CE33", X"CE2C", X"CE25", X"CE1D", X"CE16", X"CE0F", X"CE08", X"CE01", X"CDFA", X"CDF3", 
X"CDEC", X"CDE5", X"CDDE", X"CDD7", X"CDD0", X"CDC8", X"CDC1", X"CDBA", X"CDB3", X"CDAC", 
X"CDA5", X"CD9E", X"CD97", X"CD90", X"CD88", X"CD81", X"CD7A", X"CD73", X"CD6C", X"CD65", 
X"CD5E", X"CD57", X"CD50", X"CD48", X"CD41", X"CD3A", X"CD33", X"CD2C", X"CD25", X"CD1E", 
X"CD17", X"CD0F", X"CD08", X"CD01", X"CCFA", X"CCF3", X"CCEC", X"CCE5", X"CCDD", X"CCD6", 
X"CCCF", X"CCC8", X"CCC1", X"CCBA", X"CCB3", X"CCAB", X"CCA4", X"CC9D", X"CC96", X"CC8F", 
X"CC88", X"CC80", X"CC79", X"CC72", X"CC6B", X"CC64", X"CC5D", X"CC55", X"CC4E", X"CC47", 
X"CC40", X"CC39", X"CC32", X"CC2A", X"CC23", X"CC1C", X"CC15", X"CC0E", X"CC06", X"CBFF", 
X"CBF8", X"CBF1", X"CBEA", X"CBE2", X"CBDB", X"CBD4", X"CBCD", X"CBC6", X"CBBE", X"CBB7", 
X"CBB0", X"CBA9", X"CBA2", X"CB9A", X"CB93", X"CB8C", X"CB85", X"CB7E", X"CB76", X"CB6F", 
X"CB68", X"CB61", X"CB59", X"CB52", X"CB4B", X"CB44", X"CB3D", X"CB35", X"CB2E", X"CB27", 
X"CB20", X"CB18", X"CB11", X"CB0A", X"CB03", X"CAFB", X"CAF4", X"CAED", X"CAE6", X"CADE", 
X"CAD7", X"CAD0", X"CAC9", X"CAC1", X"CABA", X"CAB3", X"CAAC", X"CAA4", X"CA9D", X"CA96", 
X"CA8F", X"CA87", X"CA80", X"CA79", X"CA72", X"CA6A", X"CA63", X"CA5C", X"CA54", X"CA4D", 
X"CA46", X"CA3F", X"CA37", X"CA30", X"CA29", X"CA22", X"CA1A", X"CA13", X"CA0C", X"CA04", 
X"C9FD", X"C9F6", X"C9EE", X"C9E7", X"C9E0", X"C9D9", X"C9D1", X"C9CA", X"C9C3", X"C9BB", 
X"C9B4", X"C9AD", X"C9A5", X"C99E", X"C997", X"C990", X"C988", X"C981", X"C97A", X"C972", 
X"C96B", X"C964", X"C95C", X"C955", X"C94E", X"C946", X"C93F", X"C938", X"C930", X"C929", 
X"C922", X"C91A", X"C913", X"C90C", X"C904", X"C8FD", X"C8F6", X"C8EE", X"C8E7", X"C8E0", 
X"C8D8", X"C8D1", X"C8CA", X"C8C2", X"C8BB", X"C8B4", X"C8AC", X"C8A5", X"C89D", X"C896", 
X"C88F", X"C887", X"C880", X"C879", X"C871", X"C86A", X"C863", X"C85B", X"C854", X"C84C", 
X"C845", X"C83E", X"C836", X"C82F", X"C828", X"C820", X"C819", X"C811", X"C80A", X"C803", 
X"C7FB", X"C7F4", X"C7EC", X"C7E5", X"C7DE", X"C7D6", X"C7CF", X"C7C7", X"C7C0", X"C7B9", 
X"C7B1", X"C7AA", X"C7A2", X"C79B", X"C794", X"C78C", X"C785", X"C77D", X"C776", X"C76F", 
X"C767", X"C760", X"C758", X"C751", X"C749", X"C742", X"C73B", X"C733", X"C72C", X"C724", 
X"C71D", X"C715", X"C70E", X"C707", X"C6FF", X"C6F8", X"C6F0", X"C6E9", X"C6E1", X"C6DA", 
X"C6D3", X"C6CB", X"C6C4", X"C6BC", X"C6B5", X"C6AD", X"C6A6", X"C69E", X"C697", X"C690", 
X"C688", X"C681", X"C679", X"C672", X"C66A", X"C663", X"C65B", X"C654", X"C64C", X"C645", 
X"C63D", X"C636", X"C62E", X"C627", X"C620", X"C618", X"C611", X"C609", X"C602", X"C5FA", 
X"C5F3", X"C5EB", X"C5E4", X"C5DC", X"C5D5", X"C5CD", X"C5C6", X"C5BE", X"C5B7", X"C5AF", 
X"C5A8", X"C5A0", X"C599", X"C591", X"C58A", X"C582", X"C57B", X"C573", X"C56C", X"C564", 
X"C55D", X"C555", X"C54E", X"C546", X"C53F", X"C537", X"C530", X"C528", X"C521", X"C519", 
X"C512", X"C50A", X"C502", X"C4FB", X"C4F3", X"C4EC", X"C4E4", X"C4DD", X"C4D5", X"C4CE", 
X"C4C6", X"C4BF", X"C4B7", X"C4B0", X"C4A8", X"C4A1", X"C499", X"C491", X"C48A", X"C482", 
X"C47B", X"C473", X"C46C", X"C464", X"C45D", X"C455", X"C44D", X"C446", X"C43E", X"C437", 
X"C42F", X"C428", X"C420", X"C419", X"C411", X"C409", X"C402", X"C3FA", X"C3F3", X"C3EB", 
X"C3E4", X"C3DC", X"C3D4", X"C3CD", X"C3C5", X"C3BE", X"C3B6", X"C3AE", X"C3A7", X"C39F", 
X"C398", X"C390", X"C389", X"C381", X"C379", X"C372", X"C36A", X"C363", X"C35B", X"C353", 
X"C34C", X"C344", X"C33D", X"C335", X"C32D", X"C326", X"C31E", X"C317", X"C30F", X"C307", 
X"C300", X"C2F8", X"C2F0", X"C2E9", X"C2E1", X"C2DA", X"C2D2", X"C2CA", X"C2C3", X"C2BB", 
X"C2B3", X"C2AC", X"C2A4", X"C29D", X"C295", X"C28D", X"C286", X"C27E", X"C276", X"C26F", 
X"C267", X"C260", X"C258", X"C250", X"C249", X"C241", X"C239", X"C232", X"C22A", X"C222", 
X"C21B", X"C213", X"C20B", X"C204", X"C1FC", X"C1F4", X"C1ED", X"C1E5", X"C1DD", X"C1D6", 
X"C1CE", X"C1C6", X"C1BF", X"C1B7", X"C1AF", X"C1A8", X"C1A0", X"C198", X"C191", X"C189", 
X"C181", X"C17A", X"C172", X"C16A", X"C163", X"C15B", X"C153", X"C14C", X"C144", X"C13C", 
X"C135", X"C12D", X"C125", X"C11E", X"C116", X"C10E", X"C106", X"C0FF", X"C0F7", X"C0EF", 
X"C0E8", X"C0E0", X"C0D8", X"C0D1", X"C0C9", X"C0C1", X"C0B9", X"C0B2", X"C0AA", X"C0A2", 
X"C09B", X"C093", X"C08B", X"C083", X"C07C", X"C074", X"C06C", X"C065", X"C05D", X"C055", 
X"C04D", X"C046", X"C03E", X"C036", X"C02E", X"C027", X"C01F", X"C017", X"C00F", X"C008", 
X"C000", X"BFF8", X"BFF1", X"BFE9", X"BFE1", X"BFD9", X"BFD2", X"BFCA", X"BFC2", X"BFBA", 
X"BFB3", X"BFAB", X"BFA3", X"BF9B", X"BF94", X"BF8C", X"BF84", X"BF7C", X"BF75", X"BF6D", 
X"BF65", X"BF5D", X"BF55", X"BF4E", X"BF46", X"BF3E", X"BF36", X"BF2F", X"BF27", X"BF1F", 
X"BF17", X"BF10", X"BF08", X"BF00", X"BEF8", X"BEF0", X"BEE9", X"BEE1", X"BED9", X"BED1", 
X"BEC9", X"BEC2", X"BEBA", X"BEB2", X"BEAA", X"BEA3", X"BE9B", X"BE93", X"BE8B", X"BE83", 
X"BE7C", X"BE74", X"BE6C", X"BE64", X"BE5C", X"BE55", X"BE4D", X"BE45", X"BE3D", X"BE35", 
X"BE2D", X"BE26", X"BE1E", X"BE16", X"BE0E", X"BE06", X"BDFF", X"BDF7", X"BDEF", X"BDE7", 
X"BDDF", X"BDD8", X"BDD0", X"BDC8", X"BDC0", X"BDB8", X"BDB0", X"BDA9", X"BDA1", X"BD99", 
X"BD91", X"BD89", X"BD81", X"BD7A", X"BD72", X"BD6A", X"BD62", X"BD5A", X"BD52", X"BD4A", 
X"BD43", X"BD3B", X"BD33", X"BD2B", X"BD23", X"BD1B", X"BD14", X"BD0C", X"BD04", X"BCFC", 
X"BCF4", X"BCEC", X"BCE4", X"BCDD", X"BCD5", X"BCCD", X"BCC5", X"BCBD", X"BCB5", X"BCAD", 
X"BCA5", X"BC9E", X"BC96", X"BC8E", X"BC86", X"BC7E", X"BC76", X"BC6E", X"BC66", X"BC5F", 
X"BC57", X"BC4F", X"BC47", X"BC3F", X"BC37", X"BC2F", X"BC27", X"BC20", X"BC18", X"BC10", 
X"BC08", X"BC00", X"BBF8", X"BBF0", X"BBE8", X"BBE0", X"BBD8", X"BBD1", X"BBC9", X"BBC1", 
X"BBB9", X"BBB1", X"BBA9", X"BBA1", X"BB99", X"BB91", X"BB89", X"BB82", X"BB7A", X"BB72", 
X"BB6A", X"BB62", X"BB5A", X"BB52", X"BB4A", X"BB42", X"BB3A", X"BB32", X"BB2A", X"BB23", 
X"BB1B", X"BB13", X"BB0B", X"BB03", X"BAFB", X"BAF3", X"BAEB", X"BAE3", X"BADB", X"BAD3", 
X"BACB", X"BAC3", X"BABB", X"BAB3", X"BAAB", X"BAA4", X"BA9C", X"BA94", X"BA8C", X"BA84", 
X"BA7C", X"BA74", X"BA6C", X"BA64", X"BA5C", X"BA54", X"BA4C", X"BA44", X"BA3C", X"BA34", 
X"BA2C", X"BA24", X"BA1C", X"BA14", X"BA0C", X"BA04", X"B9FD", X"B9F5", X"B9ED", X"B9E5", 
X"B9DD", X"B9D5", X"B9CD", X"B9C5", X"B9BD", X"B9B5", X"B9AD", X"B9A5", X"B99D", X"B995", 
X"B98D", X"B985", X"B97D", X"B975", X"B96D", X"B965", X"B95D", X"B955", X"B94D", X"B945", 
X"B93D", X"B935", X"B92D", X"B925", X"B91D", X"B915", X"B90D", X"B905", X"B8FD", X"B8F5", 
X"B8ED", X"B8E5", X"B8DD", X"B8D5", X"B8CD", X"B8C5", X"B8BD", X"B8B5", X"B8AD", X"B8A5", 
X"B89D", X"B895", X"B88D", X"B885", X"B87D", X"B875", X"B86D", X"B865", X"B85D", X"B855", 
X"B84D", X"B845", X"B83D", X"B835", X"B82D", X"B825", X"B81D", X"B815", X"B80C", X"B804", 
X"B7FC", X"B7F4", X"B7EC", X"B7E4", X"B7DC", X"B7D4", X"B7CC", X"B7C4", X"B7BC", X"B7B4", 
X"B7AC", X"B7A4", X"B79C", X"B794", X"B78C", X"B784", X"B77C", X"B774", X"B76C", X"B764", 
X"B75B", X"B753", X"B74B", X"B743", X"B73B", X"B733", X"B72B", X"B723", X"B71B", X"B713", 
X"B70B", X"B703", X"B6FB", X"B6F3", X"B6EB", X"B6E3", X"B6DA", X"B6D2", X"B6CA", X"B6C2", 
X"B6BA", X"B6B2", X"B6AA", X"B6A2", X"B69A", X"B692", X"B68A", X"B682", X"B679", X"B671", 
X"B669", X"B661", X"B659", X"B651", X"B649", X"B641", X"B639", X"B631", X"B629", X"B620", 
X"B618", X"B610", X"B608", X"B600", X"B5F8", X"B5F0", X"B5E8", X"B5E0", X"B5D8", X"B5CF", 
X"B5C7", X"B5BF", X"B5B7", X"B5AF", X"B5A7", X"B59F", X"B597", X"B58F", X"B586", X"B57E", 
X"B576", X"B56E", X"B566", X"B55E", X"B556", X"B54E", X"B545", X"B53D", X"B535", X"B52D", 
X"B525", X"B51D", X"B515", X"B50D", X"B504", X"B4FC", X"B4F4", X"B4EC", X"B4E4", X"B4DC", 
X"B4D4", X"B4CB", X"B4C3", X"B4BB", X"B4B3", X"B4AB", X"B4A3", X"B49B", X"B492", X"B48A", 
X"B482", X"B47A", X"B472", X"B46A", X"B462", X"B459", X"B451", X"B449", X"B441", X"B439", 
X"B431", X"B428", X"B420", X"B418", X"B410", X"B408", X"B400", X"B3F7", X"B3EF", X"B3E7", 
X"B3DF", X"B3D7", X"B3CF", X"B3C6", X"B3BE", X"B3B6", X"B3AE", X"B3A6", X"B39E", X"B395", 
X"B38D", X"B385", X"B37D", X"B375", X"B36C", X"B364", X"B35C", X"B354", X"B34C", X"B344", 
X"B33B", X"B333", X"B32B", X"B323", X"B31B", X"B312", X"B30A", X"B302", X"B2FA", X"B2F2", 
X"B2E9", X"B2E1", X"B2D9", X"B2D1", X"B2C9", X"B2C0", X"B2B8", X"B2B0", X"B2A8", X"B2A0", 
X"B297", X"B28F", X"B287", X"B27F", X"B277", X"B26E", X"B266", X"B25E", X"B256", X"B24D", 
X"B245", X"B23D", X"B235", X"B22D", X"B224", X"B21C", X"B214", X"B20C", X"B203", X"B1FB", 
X"B1F3", X"B1EB", X"B1E3", X"B1DA", X"B1D2", X"B1CA", X"B1C2", X"B1B9", X"B1B1", X"B1A9", 
X"B1A1", X"B198", X"B190", X"B188", X"B180", X"B178", X"B16F", X"B167", X"B15F", X"B157", 
X"B14E", X"B146", X"B13E", X"B136", X"B12D", X"B125", X"B11D", X"B115", X"B10C", X"B104", 
X"B0FC", X"B0F4", X"B0EB", X"B0E3", X"B0DB", X"B0D2", X"B0CA", X"B0C2", X"B0BA", X"B0B1", 
X"B0A9", X"B0A1", X"B099", X"B090", X"B088", X"B080", X"B078", X"B06F", X"B067", X"B05F", 
X"B056", X"B04E", X"B046", X"B03E", X"B035", X"B02D", X"B025", X"B01D", X"B014", X"B00C", 
X"B004", X"AFFB", X"AFF3", X"AFEB", X"AFE3", X"AFDA", X"AFD2", X"AFCA", X"AFC1", X"AFB9", 
X"AFB1", X"AFA9", X"AFA0", X"AF98", X"AF90", X"AF87", X"AF7F", X"AF77", X"AF6E", X"AF66", 
X"AF5E", X"AF56", X"AF4D", X"AF45", X"AF3D", X"AF34", X"AF2C", X"AF24", X"AF1B", X"AF13", 
X"AF0B", X"AF02", X"AEFA", X"AEF2", X"AEEA", X"AEE1", X"AED9", X"AED1", X"AEC8", X"AEC0", 
X"AEB8", X"AEAF", X"AEA7", X"AE9F", X"AE96", X"AE8E", X"AE86", X"AE7D", X"AE75", X"AE6D", 
X"AE64", X"AE5C", X"AE54", X"AE4B", X"AE43", X"AE3B", X"AE32", X"AE2A", X"AE22", X"AE19", 
X"AE11", X"AE09", X"AE00", X"ADF8", X"ADF0", X"ADE7", X"ADDF", X"ADD7", X"ADCE", X"ADC6", 
X"ADBE", X"ADB5", X"ADAD", X"ADA5", X"AD9C", X"AD94", X"AD8C", X"AD83", X"AD7B", X"AD72", 
X"AD6A", X"AD62", X"AD59", X"AD51", X"AD49", X"AD40", X"AD38", X"AD30", X"AD27", X"AD1F", 
X"AD17", X"AD0E", X"AD06", X"ACFD", X"ACF5", X"ACED", X"ACE4", X"ACDC", X"ACD4", X"ACCB", 
X"ACC3", X"ACBA", X"ACB2", X"ACAA", X"ACA1", X"AC99", X"AC91", X"AC88", X"AC80", X"AC77", 
X"AC6F", X"AC67", X"AC5E", X"AC56", X"AC4E", X"AC45", X"AC3D", X"AC34", X"AC2C", X"AC24", 
X"AC1B", X"AC13", X"AC0A", X"AC02", X"ABFA", X"ABF1", X"ABE9", X"ABE1", X"ABD8", X"ABD0", 
X"ABC7", X"ABBF", X"ABB7", X"ABAE", X"ABA6", X"AB9D", X"AB95", X"AB8D", X"AB84", X"AB7C", 
X"AB73", X"AB6B", X"AB62", X"AB5A", X"AB52", X"AB49", X"AB41", X"AB38", X"AB30", X"AB28", 
X"AB1F", X"AB17", X"AB0E", X"AB06", X"AAFE", X"AAF5", X"AAED", X"AAE4", X"AADC", X"AAD3", 
X"AACB", X"AAC3", X"AABA", X"AAB2", X"AAA9", X"AAA1", X"AA98", X"AA90", X"AA88", X"AA7F", 
X"AA77", X"AA6E", X"AA66", X"AA5D", X"AA55", X"AA4D", X"AA44", X"AA3C", X"AA33", X"AA2B", 
X"AA22", X"AA1A", X"AA12", X"AA09", X"AA01", X"A9F8", X"A9F0", X"A9E7", X"A9DF", X"A9D6", 
X"A9CE", X"A9C6", X"A9BD", X"A9B5", X"A9AC", X"A9A4", X"A99B", X"A993", X"A98A", X"A982", 
X"A97A", X"A971", X"A969", X"A960", X"A958", X"A94F", X"A947", X"A93E", X"A936", X"A92D", 
X"A925", X"A91C", X"A914", X"A90C", X"A903", X"A8FB", X"A8F2", X"A8EA", X"A8E1", X"A8D9", 
X"A8D0", X"A8C8", X"A8BF", X"A8B7", X"A8AE", X"A8A6", X"A89D", X"A895", X"A88C", X"A884", 
X"A87C", X"A873", X"A86B", X"A862", X"A85A", X"A851", X"A849", X"A840", X"A838", X"A82F", 
X"A827", X"A81E", X"A816", X"A80D", X"A805", X"A7FC", X"A7F4", X"A7EB", X"A7E3", X"A7DA", 
X"A7D2", X"A7C9", X"A7C1", X"A7B8", X"A7B0", X"A7A7", X"A79F", X"A796", X"A78E", X"A785", 
X"A77D", X"A774", X"A76C", X"A763", X"A75B", X"A752", X"A74A", X"A741", X"A739", X"A730", 
X"A728", X"A71F", X"A717", X"A70E", X"A706", X"A6FD", X"A6F5", X"A6EC", X"A6E4", X"A6DB", 
X"A6D3", X"A6CA", X"A6C2", X"A6B9", X"A6B1", X"A6A8", X"A6A0", X"A697", X"A68F", X"A686", 
X"A67E", X"A675", X"A66C", X"A664", X"A65B", X"A653", X"A64A", X"A642", X"A639", X"A631", 
X"A628", X"A620", X"A617", X"A60F", X"A606", X"A5FE", X"A5F5", X"A5ED", X"A5E4", X"A5DB", 
X"A5D3", X"A5CA", X"A5C2", X"A5B9", X"A5B1", X"A5A8", X"A5A0", X"A597", X"A58F", X"A586", 
X"A57E", X"A575", X"A56C", X"A564", X"A55B", X"A553", X"A54A", X"A542", X"A539", X"A531", 
X"A528", X"A51F", X"A517", X"A50E", X"A506", X"A4FD", X"A4F5", X"A4EC", X"A4E4", X"A4DB", 
X"A4D3", X"A4CA", X"A4C1", X"A4B9", X"A4B0", X"A4A8", X"A49F", X"A497", X"A48E", X"A485", 
X"A47D", X"A474", X"A46C", X"A463", X"A45B", X"A452", X"A449", X"A441", X"A438", X"A430", 
X"A427", X"A41F", X"A416", X"A40D", X"A405", X"A3FC", X"A3F4", X"A3EB", X"A3E3", X"A3DA", 
X"A3D1", X"A3C9", X"A3C0", X"A3B8", X"A3AF", X"A3A7", X"A39E", X"A395", X"A38D", X"A384", 
X"A37C", X"A373", X"A36A", X"A362", X"A359", X"A351", X"A348", X"A33F", X"A337", X"A32E", 
X"A326", X"A31D", X"A315", X"A30C", X"A303", X"A2FB", X"A2F2", X"A2EA", X"A2E1", X"A2D8", 
X"A2D0", X"A2C7", X"A2BF", X"A2B6", X"A2AD", X"A2A5", X"A29C", X"A294", X"A28B", X"A282", 
X"A27A", X"A271", X"A269", X"A260", X"A257", X"A24F", X"A246", X"A23D", X"A235", X"A22C", 
X"A224", X"A21B", X"A212", X"A20A", X"A201", X"A1F9", X"A1F0", X"A1E7", X"A1DF", X"A1D6", 
X"A1CD", X"A1C5", X"A1BC", X"A1B4", X"A1AB", X"A1A2", X"A19A", X"A191", X"A189", X"A180", 
X"A177", X"A16F", X"A166", X"A15D", X"A155", X"A14C", X"A144", X"A13B", X"A132", X"A12A", 
X"A121", X"A118", X"A110", X"A107", X"A0FE", X"A0F6", X"A0ED", X"A0E5", X"A0DC", X"A0D3", 
X"A0CB", X"A0C2", X"A0B9", X"A0B1", X"A0A8", X"A09F", X"A097", X"A08E", X"A086", X"A07D", 
X"A074", X"A06C", X"A063", X"A05A", X"A052", X"A049", X"A040", X"A038", X"A02F", X"A026", 
X"A01E", X"A015", X"A00C", X"A004", X"9FFB", X"9FF2", X"9FEA", X"9FE1", X"9FD9", X"9FD0", 
X"9FC7", X"9FBF", X"9FB6", X"9FAD", X"9FA5", X"9F9C", X"9F93", X"9F8B", X"9F82", X"9F79", 
X"9F71", X"9F68", X"9F5F", X"9F57", X"9F4E", X"9F45", X"9F3D", X"9F34", X"9F2B", X"9F23", 
X"9F1A", X"9F11", X"9F09", X"9F00", X"9EF7", X"9EEF", X"9EE6", X"9EDD", X"9ED5", X"9ECC", 
X"9EC3", X"9EBB", X"9EB2", X"9EA9", X"9EA1", X"9E98", X"9E8F", X"9E87", X"9E7E", X"9E75", 
X"9E6C", X"9E64", X"9E5B", X"9E52", X"9E4A", X"9E41", X"9E38", X"9E30", X"9E27", X"9E1E", 
X"9E16", X"9E0D", X"9E04", X"9DFC", X"9DF3", X"9DEA", X"9DE2", X"9DD9", X"9DD0", X"9DC7", 
X"9DBF", X"9DB6", X"9DAD", X"9DA5", X"9D9C", X"9D93", X"9D8B", X"9D82", X"9D79", X"9D71", 
X"9D68", X"9D5F", X"9D56", X"9D4E", X"9D45", X"9D3C", X"9D34", X"9D2B", X"9D22", X"9D1A", 
X"9D11", X"9D08", X"9CFF", X"9CF7", X"9CEE", X"9CE5", X"9CDD", X"9CD4", X"9CCB", X"9CC2", 
X"9CBA", X"9CB1", X"9CA8", X"9CA0", X"9C97", X"9C8E", X"9C86", X"9C7D", X"9C74", X"9C6B", 
X"9C63", X"9C5A", X"9C51", X"9C49", X"9C40", X"9C37", X"9C2E", X"9C26", X"9C1D", X"9C14", 
X"9C0C", X"9C03", X"9BFA", X"9BF1", X"9BE9", X"9BE0", X"9BD7", X"9BCE", X"9BC6", X"9BBD", 
X"9BB4", X"9BAC", X"9BA3", X"9B9A", X"9B91", X"9B89", X"9B80", X"9B77", X"9B6E", X"9B66", 
X"9B5D", X"9B54", X"9B4C", X"9B43", X"9B3A", X"9B31", X"9B29", X"9B20", X"9B17", X"9B0E", 
X"9B06", X"9AFD", X"9AF4", X"9AEB", X"9AE3", X"9ADA", X"9AD1", X"9AC9", X"9AC0", X"9AB7", 
X"9AAE", X"9AA6", X"9A9D", X"9A94", X"9A8B", X"9A83", X"9A7A", X"9A71", X"9A68", X"9A60", 
X"9A57", X"9A4E", X"9A45", X"9A3D", X"9A34", X"9A2B", X"9A22", X"9A1A", X"9A11", X"9A08", 
X"99FF", X"99F7", X"99EE", X"99E5", X"99DC", X"99D4", X"99CB", X"99C2", X"99B9", X"99B1", 
X"99A8", X"999F", X"9996", X"998E", X"9985", X"997C", X"9973", X"996B", X"9962", X"9959", 
X"9950", X"9948", X"993F", X"9936", X"992D", X"9925", X"991C", X"9913", X"990A", X"9901", 
X"98F9", X"98F0", X"98E7", X"98DE", X"98D6", X"98CD", X"98C4", X"98BB", X"98B3", X"98AA", 
X"98A1", X"9898", X"9890", X"9887", X"987E", X"9875", X"986C", X"9864", X"985B", X"9852", 
X"9849", X"9841", X"9838", X"982F", X"9826", X"981D", X"9815", X"980C", X"9803", X"97FA", 
X"97F2", X"97E9", X"97E0", X"97D7", X"97CE", X"97C6", X"97BD", X"97B4", X"97AB", X"97A3", 
X"979A", X"9791", X"9788", X"977F", X"9777", X"976E", X"9765", X"975C", X"9753", X"974B", 
X"9742", X"9739", X"9730", X"9728", X"971F", X"9716", X"970D", X"9704", X"96FC", X"96F3", 
X"96EA", X"96E1", X"96D8", X"96D0", X"96C7", X"96BE", X"96B5", X"96AC", X"96A4", X"969B", 
X"9692", X"9689", X"9680", X"9678", X"966F", X"9666", X"965D", X"9655", X"964C", X"9643", 
X"963A", X"9631", X"9629", X"9620", X"9617", X"960E", X"9605", X"95FC", X"95F4", X"95EB", 
X"95E2", X"95D9", X"95D0", X"95C8", X"95BF", X"95B6", X"95AD", X"95A4", X"959C", X"9593", 
X"958A", X"9581", X"9578", X"9570", X"9567", X"955E", X"9555", X"954C", X"9544", X"953B", 
X"9532", X"9529", X"9520", X"9517", X"950F", X"9506", X"94FD", X"94F4", X"94EB", X"94E3", 
X"94DA", X"94D1", X"94C8", X"94BF", X"94B6", X"94AE", X"94A5", X"949C", X"9493", X"948A", 
X"9482", X"9479", X"9470", X"9467", X"945E", X"9455", X"944D", X"9444", X"943B", X"9432", 
X"9429", X"9421", X"9418", X"940F", X"9406", X"93FD", X"93F4", X"93EC", X"93E3", X"93DA", 
X"93D1", X"93C8", X"93BF", X"93B7", X"93AE", X"93A5", X"939C", X"9393", X"938A", X"9382", 
X"9379", X"9370", X"9367", X"935E", X"9355", X"934D", X"9344", X"933B", X"9332", X"9329", 
X"9320", X"9318", X"930F", X"9306", X"92FD", X"92F4", X"92EB", X"92E3", X"92DA", X"92D1", 
X"92C8", X"92BF", X"92B6", X"92AE", X"92A5", X"929C", X"9293", X"928A", X"9281", X"9278", 
X"9270", X"9267", X"925E", X"9255", X"924C", X"9243", X"923B", X"9232", X"9229", X"9220", 
X"9217", X"920E", X"9206", X"91FD", X"91F4", X"91EB", X"91E2", X"91D9", X"91D0", X"91C8", 
X"91BF", X"91B6", X"91AD", X"91A4", X"919B", X"9192", X"918A", X"9181", X"9178", X"916F", 
X"9166", X"915D", X"9155", X"914C", X"9143", X"913A", X"9131", X"9128", X"911F", X"9117", 
X"910E", X"9105", X"90FC", X"90F3", X"90EA", X"90E1", X"90D9", X"90D0", X"90C7", X"90BE", 
X"90B5", X"90AC", X"90A3", X"909B", X"9092", X"9089", X"9080", X"9077", X"906E", X"9065", 
X"905C", X"9054", X"904B", X"9042", X"9039", X"9030", X"9027", X"901E", X"9016", X"900D", 
X"9004", X"8FFB", X"8FF2", X"8FE9", X"8FE0", X"8FD7", X"8FCF", X"8FC6", X"8FBD", X"8FB4", 
X"8FAB", X"8FA2", X"8F99", X"8F91", X"8F88", X"8F7F", X"8F76", X"8F6D", X"8F64", X"8F5B", 
X"8F52", X"8F4A", X"8F41", X"8F38", X"8F2F", X"8F26", X"8F1D", X"8F14", X"8F0B", X"8F03", 
X"8EFA", X"8EF1", X"8EE8", X"8EDF", X"8ED6", X"8ECD", X"8EC4", X"8EBC", X"8EB3", X"8EAA", 
X"8EA1", X"8E98", X"8E8F", X"8E86", X"8E7D", X"8E75", X"8E6C", X"8E63", X"8E5A", X"8E51", 
X"8E48", X"8E3F", X"8E36", X"8E2E", X"8E25", X"8E1C", X"8E13", X"8E0A", X"8E01", X"8DF8", 
X"8DEF", X"8DE6", X"8DDE", X"8DD5", X"8DCC", X"8DC3", X"8DBA", X"8DB1", X"8DA8", X"8D9F", 
X"8D97", X"8D8E", X"8D85", X"8D7C", X"8D73", X"8D6A", X"8D61", X"8D58", X"8D4F", X"8D47", 
X"8D3E", X"8D35", X"8D2C", X"8D23", X"8D1A", X"8D11", X"8D08", X"8CFF", X"8CF7", X"8CEE", 
X"8CE5", X"8CDC", X"8CD3", X"8CCA", X"8CC1", X"8CB8", X"8CAF", X"8CA7", X"8C9E", X"8C95", 
X"8C8C", X"8C83", X"8C7A", X"8C71", X"8C68", X"8C5F", X"8C56", X"8C4E", X"8C45", X"8C3C", 
X"8C33", X"8C2A", X"8C21", X"8C18", X"8C0F", X"8C06", X"8BFE", X"8BF5", X"8BEC", X"8BE3", 
X"8BDA", X"8BD1", X"8BC8", X"8BBF", X"8BB6", X"8BAD", X"8BA5", X"8B9C", X"8B93", X"8B8A", 
X"8B81", X"8B78", X"8B6F", X"8B66", X"8B5D", X"8B54", X"8B4C", X"8B43", X"8B3A", X"8B31", 
X"8B28", X"8B1F", X"8B16", X"8B0D", X"8B04", X"8AFB", X"8AF3", X"8AEA", X"8AE1", X"8AD8", 
X"8ACF", X"8AC6", X"8ABD", X"8AB4", X"8AAB", X"8AA2", X"8A99", X"8A91", X"8A88", X"8A7F", 
X"8A76", X"8A6D", X"8A64", X"8A5B", X"8A52", X"8A49", X"8A40", X"8A37", X"8A2F", X"8A26", 
X"8A1D", X"8A14", X"8A0B", X"8A02", X"89F9", X"89F0", X"89E7", X"89DE", X"89D5", X"89CD", 
X"89C4", X"89BB", X"89B2", X"89A9", X"89A0", X"8997", X"898E", X"8985", X"897C", X"8973", 
X"896B", X"8962", X"8959", X"8950", X"8947", X"893E", X"8935", X"892C", X"8923", X"891A", 
X"8911", X"8909", X"8900", X"88F7", X"88EE", X"88E5", X"88DC", X"88D3", X"88CA", X"88C1", 
X"88B8", X"88AF", X"88A6", X"889E", X"8895", X"888C", X"8883", X"887A", X"8871", X"8868", 
X"885F", X"8856", X"884D", X"8844", X"883B", X"8833", X"882A", X"8821", X"8818", X"880F", 
X"8806", X"87FD", X"87F4", X"87EB", X"87E2", X"87D9", X"87D0", X"87C8", X"87BF", X"87B6", 
X"87AD", X"87A4", X"879B", X"8792", X"8789", X"8780", X"8777", X"876E", X"8765", X"875C", 
X"8754", X"874B", X"8742", X"8739", X"8730", X"8727", X"871E", X"8715", X"870C", X"8703", 
X"86FA", X"86F1", X"86E8", X"86E0", X"86D7", X"86CE", X"86C5", X"86BC", X"86B3", X"86AA", 
X"86A1", X"8698", X"868F", X"8686", X"867D", X"8674", X"866C", X"8663", X"865A", X"8651", 
X"8648", X"863F", X"8636", X"862D", X"8624", X"861B", X"8612", X"8609", X"8600", X"85F8", 
X"85EF", X"85E6", X"85DD", X"85D4", X"85CB", X"85C2", X"85B9", X"85B0", X"85A7", X"859E", 
X"8595", X"858C", X"8583", X"857B", X"8572", X"8569", X"8560", X"8557", X"854E", X"8545", 
X"853C", X"8533", X"852A", X"8521", X"8518", X"850F", X"8506", X"84FE", X"84F5", X"84EC", 
X"84E3", X"84DA", X"84D1", X"84C8", X"84BF", X"84B6", X"84AD", X"84A4", X"849B", X"8492", 
X"8489", X"8481", X"8478", X"846F", X"8466", X"845D", X"8454", X"844B", X"8442", X"8439", 
X"8430", X"8427", X"841E", X"8415", X"840C", X"8403", X"83FB", X"83F2", X"83E9", X"83E0", 
X"83D7", X"83CE", X"83C5", X"83BC", X"83B3", X"83AA", X"83A1", X"8398", X"838F", X"8386", 
X"837D", X"8375", X"836C", X"8363", X"835A", X"8351", X"8348", X"833F", X"8336", X"832D", 
X"8324", X"831B", X"8312", X"8309", X"8300", X"82F7", X"82EF", X"82E6", X"82DD", X"82D4", 
X"82CB", X"82C2", X"82B9", X"82B0", X"82A7", X"829E", X"8295", X"828C", X"8283", X"827A", 
X"8271", X"8269", X"8260", X"8257", X"824E", X"8245", X"823C", X"8233", X"822A", X"8221", 
X"8218", X"820F", X"8206", X"81FD", X"81F4", X"81EB", X"81E3", X"81DA", X"81D1", X"81C8", 
X"81BF", X"81B6", X"81AD", X"81A4", X"819B", X"8192", X"8189", X"8180", X"8177", X"816E", 
X"8165", X"815D", X"8154", X"814B", X"8142", X"8139", X"8130", X"8127", X"811E", X"8115", 
X"810C", X"8103", X"80FA", X"80F1", X"80E8", X"80DF", X"80D6", X"80CE", X"80C5", X"80BC", 
X"80B3", X"80AA", X"80A1", X"8098", X"808F", X"8086", X"807D", X"8074", X"806B", X"8062", 
X"8059", X"8050", X"8047", X"803F", X"8036", X"802D", X"8024", X"801B", X"8012", X"8009", 
X"0000", X"0009", X"0012", X"001B", X"0024", X"002D", X"0036", X"003F", X"0047", X"0050", 
X"0059", X"0062", X"006B", X"0074", X"007D", X"0086", X"008F", X"0098", X"00A1", X"00AA", 
X"00B3", X"00BC", X"00C5", X"00CE", X"00D6", X"00DF", X"00E8", X"00F1", X"00FA", X"0103", 
X"010C", X"0115", X"011E", X"0127", X"0130", X"0139", X"0142", X"014B", X"0154", X"015D", 
X"0165", X"016E", X"0177", X"0180", X"0189", X"0192", X"019B", X"01A4", X"01AD", X"01B6", 
X"01BF", X"01C8", X"01D1", X"01DA", X"01E3", X"01EB", X"01F4", X"01FD", X"0206", X"020F", 
X"0218", X"0221", X"022A", X"0233", X"023C", X"0245", X"024E", X"0257", X"0260", X"0269", 
X"0271", X"027A", X"0283", X"028C", X"0295", X"029E", X"02A7", X"02B0", X"02B9", X"02C2", 
X"02CB", X"02D4", X"02DD", X"02E6", X"02EF", X"02F7", X"0300", X"0309", X"0312", X"031B", 
X"0324", X"032D", X"0336", X"033F", X"0348", X"0351", X"035A", X"0363", X"036C", X"0375", 
X"037D", X"0386", X"038F", X"0398", X"03A1", X"03AA", X"03B3", X"03BC", X"03C5", X"03CE", 
X"03D7", X"03E0", X"03E9", X"03F2", X"03FB", X"0403", X"040C", X"0415", X"041E", X"0427", 
X"0430", X"0439", X"0442", X"044B", X"0454", X"045D", X"0466", X"046F", X"0478", X"0481", 
X"0489", X"0492", X"049B", X"04A4", X"04AD", X"04B6", X"04BF", X"04C8", X"04D1", X"04DA", 
X"04E3", X"04EC", X"04F5", X"04FE", X"0506", X"050F", X"0518", X"0521", X"052A", X"0533", 
X"053C", X"0545", X"054E", X"0557", X"0560", X"0569", X"0572", X"057B", X"0583", X"058C", 
X"0595", X"059E", X"05A7", X"05B0", X"05B9", X"05C2", X"05CB", X"05D4", X"05DD", X"05E6", 
X"05EF", X"05F8", X"0600", X"0609", X"0612", X"061B", X"0624", X"062D", X"0636", X"063F", 
X"0648", X"0651", X"065A", X"0663", X"066C", X"0674", X"067D", X"0686", X"068F", X"0698", 
X"06A1", X"06AA", X"06B3", X"06BC", X"06C5", X"06CE", X"06D7", X"06E0", X"06E8", X"06F1", 
X"06FA", X"0703", X"070C", X"0715", X"071E", X"0727", X"0730", X"0739", X"0742", X"074B", 
X"0754", X"075C", X"0765", X"076E", X"0777", X"0780", X"0789", X"0792", X"079B", X"07A4", 
X"07AD", X"07B6", X"07BF", X"07C8", X"07D0", X"07D9", X"07E2", X"07EB", X"07F4", X"07FD", 
X"0806", X"080F", X"0818", X"0821", X"082A", X"0833", X"083B", X"0844", X"084D", X"0856", 
X"085F", X"0868", X"0871", X"087A", X"0883", X"088C", X"0895", X"089E", X"08A6", X"08AF", 
X"08B8", X"08C1", X"08CA", X"08D3", X"08DC", X"08E5", X"08EE", X"08F7", X"0900", X"0909", 
X"0911", X"091A", X"0923", X"092C", X"0935", X"093E", X"0947", X"0950", X"0959", X"0962", 
X"096B", X"0973", X"097C", X"0985", X"098E", X"0997", X"09A0", X"09A9", X"09B2", X"09BB", 
X"09C4", X"09CD", X"09D5", X"09DE", X"09E7", X"09F0", X"09F9", X"0A02", X"0A0B", X"0A14", 
X"0A1D", X"0A26", X"0A2F", X"0A37", X"0A40", X"0A49", X"0A52", X"0A5B", X"0A64", X"0A6D", 
X"0A76", X"0A7F", X"0A88", X"0A91", X"0A99", X"0AA2", X"0AAB", X"0AB4", X"0ABD", X"0AC6", 
X"0ACF", X"0AD8", X"0AE1", X"0AEA", X"0AF3", X"0AFB", X"0B04", X"0B0D", X"0B16", X"0B1F", 
X"0B28", X"0B31", X"0B3A", X"0B43", X"0B4C", X"0B54", X"0B5D", X"0B66", X"0B6F", X"0B78", 
X"0B81", X"0B8A", X"0B93", X"0B9C", X"0BA5", X"0BAD", X"0BB6", X"0BBF", X"0BC8", X"0BD1", 
X"0BDA", X"0BE3", X"0BEC", X"0BF5", X"0BFE", X"0C06", X"0C0F", X"0C18", X"0C21", X"0C2A", 
X"0C33", X"0C3C", X"0C45", X"0C4E", X"0C56", X"0C5F", X"0C68", X"0C71", X"0C7A", X"0C83", 
X"0C8C", X"0C95", X"0C9E", X"0CA7", X"0CAF", X"0CB8", X"0CC1", X"0CCA", X"0CD3", X"0CDC", 
X"0CE5", X"0CEE", X"0CF7", X"0CFF", X"0D08", X"0D11", X"0D1A", X"0D23", X"0D2C", X"0D35", 
X"0D3E", X"0D47", X"0D4F", X"0D58", X"0D61", X"0D6A", X"0D73", X"0D7C", X"0D85", X"0D8E", 
X"0D97", X"0D9F", X"0DA8", X"0DB1", X"0DBA", X"0DC3", X"0DCC", X"0DD5", X"0DDE", X"0DE6", 
X"0DEF", X"0DF8", X"0E01", X"0E0A", X"0E13", X"0E1C", X"0E25", X"0E2E", X"0E36", X"0E3F", 
X"0E48", X"0E51", X"0E5A", X"0E63", X"0E6C", X"0E75", X"0E7D", X"0E86", X"0E8F", X"0E98", 
X"0EA1", X"0EAA", X"0EB3", X"0EBC", X"0EC4", X"0ECD", X"0ED6", X"0EDF", X"0EE8", X"0EF1", 
X"0EFA", X"0F03", X"0F0B", X"0F14", X"0F1D", X"0F26", X"0F2F", X"0F38", X"0F41", X"0F4A", 
X"0F52", X"0F5B", X"0F64", X"0F6D", X"0F76", X"0F7F", X"0F88", X"0F91", X"0F99", X"0FA2", 
X"0FAB", X"0FB4", X"0FBD", X"0FC6", X"0FCF", X"0FD7", X"0FE0", X"0FE9", X"0FF2", X"0FFB", 
X"1004", X"100D", X"1016", X"101E", X"1027", X"1030", X"1039", X"1042", X"104B", X"1054", 
X"105C", X"1065", X"106E", X"1077", X"1080", X"1089", X"1092", X"109B", X"10A3", X"10AC", 
X"10B5", X"10BE", X"10C7", X"10D0", X"10D9", X"10E1", X"10EA", X"10F3", X"10FC", X"1105", 
X"110E", X"1117", X"111F", X"1128", X"1131", X"113A", X"1143", X"114C", X"1155", X"115D", 
X"1166", X"116F", X"1178", X"1181", X"118A", X"1192", X"119B", X"11A4", X"11AD", X"11B6", 
X"11BF", X"11C8", X"11D0", X"11D9", X"11E2", X"11EB", X"11F4", X"11FD", X"1206", X"120E", 
X"1217", X"1220", X"1229", X"1232", X"123B", X"1243", X"124C", X"1255", X"125E", X"1267", 
X"1270", X"1278", X"1281", X"128A", X"1293", X"129C", X"12A5", X"12AE", X"12B6", X"12BF", 
X"12C8", X"12D1", X"12DA", X"12E3", X"12EB", X"12F4", X"12FD", X"1306", X"130F", X"1318", 
X"1320", X"1329", X"1332", X"133B", X"1344", X"134D", X"1355", X"135E", X"1367", X"1370", 
X"1379", X"1382", X"138A", X"1393", X"139C", X"13A5", X"13AE", X"13B7", X"13BF", X"13C8", 
X"13D1", X"13DA", X"13E3", X"13EC", X"13F4", X"13FD", X"1406", X"140F", X"1418", X"1421", 
X"1429", X"1432", X"143B", X"1444", X"144D", X"1455", X"145E", X"1467", X"1470", X"1479", 
X"1482", X"148A", X"1493", X"149C", X"14A5", X"14AE", X"14B6", X"14BF", X"14C8", X"14D1", 
X"14DA", X"14E3", X"14EB", X"14F4", X"14FD", X"1506", X"150F", X"1517", X"1520", X"1529", 
X"1532", X"153B", X"1544", X"154C", X"1555", X"155E", X"1567", X"1570", X"1578", X"1581", 
X"158A", X"1593", X"159C", X"15A4", X"15AD", X"15B6", X"15BF", X"15C8", X"15D0", X"15D9", 
X"15E2", X"15EB", X"15F4", X"15FC", X"1605", X"160E", X"1617", X"1620", X"1629", X"1631", 
X"163A", X"1643", X"164C", X"1655", X"165D", X"1666", X"166F", X"1678", X"1680", X"1689", 
X"1692", X"169B", X"16A4", X"16AC", X"16B5", X"16BE", X"16C7", X"16D0", X"16D8", X"16E1", 
X"16EA", X"16F3", X"16FC", X"1704", X"170D", X"1716", X"171F", X"1728", X"1730", X"1739", 
X"1742", X"174B", X"1753", X"175C", X"1765", X"176E", X"1777", X"177F", X"1788", X"1791", 
X"179A", X"17A3", X"17AB", X"17B4", X"17BD", X"17C6", X"17CE", X"17D7", X"17E0", X"17E9", 
X"17F2", X"17FA", X"1803", X"180C", X"1815", X"181D", X"1826", X"182F", X"1838", X"1841", 
X"1849", X"1852", X"185B", X"1864", X"186C", X"1875", X"187E", X"1887", X"1890", X"1898", 
X"18A1", X"18AA", X"18B3", X"18BB", X"18C4", X"18CD", X"18D6", X"18DE", X"18E7", X"18F0", 
X"18F9", X"1901", X"190A", X"1913", X"191C", X"1925", X"192D", X"1936", X"193F", X"1948", 
X"1950", X"1959", X"1962", X"196B", X"1973", X"197C", X"1985", X"198E", X"1996", X"199F", 
X"19A8", X"19B1", X"19B9", X"19C2", X"19CB", X"19D4", X"19DC", X"19E5", X"19EE", X"19F7", 
X"19FF", X"1A08", X"1A11", X"1A1A", X"1A22", X"1A2B", X"1A34", X"1A3D", X"1A45", X"1A4E", 
X"1A57", X"1A60", X"1A68", X"1A71", X"1A7A", X"1A83", X"1A8B", X"1A94", X"1A9D", X"1AA6", 
X"1AAE", X"1AB7", X"1AC0", X"1AC9", X"1AD1", X"1ADA", X"1AE3", X"1AEB", X"1AF4", X"1AFD", 
X"1B06", X"1B0E", X"1B17", X"1B20", X"1B29", X"1B31", X"1B3A", X"1B43", X"1B4C", X"1B54", 
X"1B5D", X"1B66", X"1B6E", X"1B77", X"1B80", X"1B89", X"1B91", X"1B9A", X"1BA3", X"1BAC", 
X"1BB4", X"1BBD", X"1BC6", X"1BCE", X"1BD7", X"1BE0", X"1BE9", X"1BF1", X"1BFA", X"1C03", 
X"1C0C", X"1C14", X"1C1D", X"1C26", X"1C2E", X"1C37", X"1C40", X"1C49", X"1C51", X"1C5A", 
X"1C63", X"1C6B", X"1C74", X"1C7D", X"1C86", X"1C8E", X"1C97", X"1CA0", X"1CA8", X"1CB1", 
X"1CBA", X"1CC2", X"1CCB", X"1CD4", X"1CDD", X"1CE5", X"1CEE", X"1CF7", X"1CFF", X"1D08", 
X"1D11", X"1D1A", X"1D22", X"1D2B", X"1D34", X"1D3C", X"1D45", X"1D4E", X"1D56", X"1D5F", 
X"1D68", X"1D71", X"1D79", X"1D82", X"1D8B", X"1D93", X"1D9C", X"1DA5", X"1DAD", X"1DB6", 
X"1DBF", X"1DC7", X"1DD0", X"1DD9", X"1DE2", X"1DEA", X"1DF3", X"1DFC", X"1E04", X"1E0D", 
X"1E16", X"1E1E", X"1E27", X"1E30", X"1E38", X"1E41", X"1E4A", X"1E52", X"1E5B", X"1E64", 
X"1E6C", X"1E75", X"1E7E", X"1E87", X"1E8F", X"1E98", X"1EA1", X"1EA9", X"1EB2", X"1EBB", 
X"1EC3", X"1ECC", X"1ED5", X"1EDD", X"1EE6", X"1EEF", X"1EF7", X"1F00", X"1F09", X"1F11", 
X"1F1A", X"1F23", X"1F2B", X"1F34", X"1F3D", X"1F45", X"1F4E", X"1F57", X"1F5F", X"1F68", 
X"1F71", X"1F79", X"1F82", X"1F8B", X"1F93", X"1F9C", X"1FA5", X"1FAD", X"1FB6", X"1FBF", 
X"1FC7", X"1FD0", X"1FD9", X"1FE1", X"1FEA", X"1FF2", X"1FFB", X"2004", X"200C", X"2015", 
X"201E", X"2026", X"202F", X"2038", X"2040", X"2049", X"2052", X"205A", X"2063", X"206C", 
X"2074", X"207D", X"2086", X"208E", X"2097", X"209F", X"20A8", X"20B1", X"20B9", X"20C2", 
X"20CB", X"20D3", X"20DC", X"20E5", X"20ED", X"20F6", X"20FE", X"2107", X"2110", X"2118", 
X"2121", X"212A", X"2132", X"213B", X"2144", X"214C", X"2155", X"215D", X"2166", X"216F", 
X"2177", X"2180", X"2189", X"2191", X"219A", X"21A2", X"21AB", X"21B4", X"21BC", X"21C5", 
X"21CD", X"21D6", X"21DF", X"21E7", X"21F0", X"21F9", X"2201", X"220A", X"2212", X"221B", 
X"2224", X"222C", X"2235", X"223D", X"2246", X"224F", X"2257", X"2260", X"2269", X"2271", 
X"227A", X"2282", X"228B", X"2294", X"229C", X"22A5", X"22AD", X"22B6", X"22BF", X"22C7", 
X"22D0", X"22D8", X"22E1", X"22EA", X"22F2", X"22FB", X"2303", X"230C", X"2315", X"231D", 
X"2326", X"232E", X"2337", X"233F", X"2348", X"2351", X"2359", X"2362", X"236A", X"2373", 
X"237C", X"2384", X"238D", X"2395", X"239E", X"23A7", X"23AF", X"23B8", X"23C0", X"23C9", 
X"23D1", X"23DA", X"23E3", X"23EB", X"23F4", X"23FC", X"2405", X"240D", X"2416", X"241F", 
X"2427", X"2430", X"2438", X"2441", X"2449", X"2452", X"245B", X"2463", X"246C", X"2474", 
X"247D", X"2485", X"248E", X"2497", X"249F", X"24A8", X"24B0", X"24B9", X"24C1", X"24CA", 
X"24D3", X"24DB", X"24E4", X"24EC", X"24F5", X"24FD", X"2506", X"250E", X"2517", X"251F", 
X"2528", X"2531", X"2539", X"2542", X"254A", X"2553", X"255B", X"2564", X"256C", X"2575", 
X"257E", X"2586", X"258F", X"2597", X"25A0", X"25A8", X"25B1", X"25B9", X"25C2", X"25CA", 
X"25D3", X"25DB", X"25E4", X"25ED", X"25F5", X"25FE", X"2606", X"260F", X"2617", X"2620", 
X"2628", X"2631", X"2639", X"2642", X"264A", X"2653", X"265B", X"2664", X"266C", X"2675", 
X"267E", X"2686", X"268F", X"2697", X"26A0", X"26A8", X"26B1", X"26B9", X"26C2", X"26CA", 
X"26D3", X"26DB", X"26E4", X"26EC", X"26F5", X"26FD", X"2706", X"270E", X"2717", X"271F", 
X"2728", X"2730", X"2739", X"2741", X"274A", X"2752", X"275B", X"2763", X"276C", X"2774", 
X"277D", X"2785", X"278E", X"2796", X"279F", X"27A7", X"27B0", X"27B8", X"27C1", X"27C9", 
X"27D2", X"27DA", X"27E3", X"27EB", X"27F4", X"27FC", X"2805", X"280D", X"2816", X"281E", 
X"2827", X"282F", X"2838", X"2840", X"2849", X"2851", X"285A", X"2862", X"286B", X"2873", 
X"287C", X"2884", X"288C", X"2895", X"289D", X"28A6", X"28AE", X"28B7", X"28BF", X"28C8", 
X"28D0", X"28D9", X"28E1", X"28EA", X"28F2", X"28FB", X"2903", X"290C", X"2914", X"291C", 
X"2925", X"292D", X"2936", X"293E", X"2947", X"294F", X"2958", X"2960", X"2969", X"2971", 
X"297A", X"2982", X"298A", X"2993", X"299B", X"29A4", X"29AC", X"29B5", X"29BD", X"29C6", 
X"29CE", X"29D6", X"29DF", X"29E7", X"29F0", X"29F8", X"2A01", X"2A09", X"2A12", X"2A1A", 
X"2A22", X"2A2B", X"2A33", X"2A3C", X"2A44", X"2A4D", X"2A55", X"2A5D", X"2A66", X"2A6E", 
X"2A77", X"2A7F", X"2A88", X"2A90", X"2A98", X"2AA1", X"2AA9", X"2AB2", X"2ABA", X"2AC3", 
X"2ACB", X"2AD3", X"2ADC", X"2AE4", X"2AED", X"2AF5", X"2AFE", X"2B06", X"2B0E", X"2B17", 
X"2B1F", X"2B28", X"2B30", X"2B38", X"2B41", X"2B49", X"2B52", X"2B5A", X"2B62", X"2B6B", 
X"2B73", X"2B7C", X"2B84", X"2B8D", X"2B95", X"2B9D", X"2BA6", X"2BAE", X"2BB7", X"2BBF", 
X"2BC7", X"2BD0", X"2BD8", X"2BE1", X"2BE9", X"2BF1", X"2BFA", X"2C02", X"2C0A", X"2C13", 
X"2C1B", X"2C24", X"2C2C", X"2C34", X"2C3D", X"2C45", X"2C4E", X"2C56", X"2C5E", X"2C67", 
X"2C6F", X"2C77", X"2C80", X"2C88", X"2C91", X"2C99", X"2CA1", X"2CAA", X"2CB2", X"2CBA", 
X"2CC3", X"2CCB", X"2CD4", X"2CDC", X"2CE4", X"2CED", X"2CF5", X"2CFD", X"2D06", X"2D0E", 
X"2D17", X"2D1F", X"2D27", X"2D30", X"2D38", X"2D40", X"2D49", X"2D51", X"2D59", X"2D62", 
X"2D6A", X"2D72", X"2D7B", X"2D83", X"2D8C", X"2D94", X"2D9C", X"2DA5", X"2DAD", X"2DB5", 
X"2DBE", X"2DC6", X"2DCE", X"2DD7", X"2DDF", X"2DE7", X"2DF0", X"2DF8", X"2E00", X"2E09", 
X"2E11", X"2E19", X"2E22", X"2E2A", X"2E32", X"2E3B", X"2E43", X"2E4B", X"2E54", X"2E5C", 
X"2E64", X"2E6D", X"2E75", X"2E7D", X"2E86", X"2E8E", X"2E96", X"2E9F", X"2EA7", X"2EAF", 
X"2EB8", X"2EC0", X"2EC8", X"2ED1", X"2ED9", X"2EE1", X"2EEA", X"2EF2", X"2EFA", X"2F02", 
X"2F0B", X"2F13", X"2F1B", X"2F24", X"2F2C", X"2F34", X"2F3D", X"2F45", X"2F4D", X"2F56", 
X"2F5E", X"2F66", X"2F6E", X"2F77", X"2F7F", X"2F87", X"2F90", X"2F98", X"2FA0", X"2FA9", 
X"2FB1", X"2FB9", X"2FC1", X"2FCA", X"2FD2", X"2FDA", X"2FE3", X"2FEB", X"2FF3", X"2FFB", 
X"3004", X"300C", X"3014", X"301D", X"3025", X"302D", X"3035", X"303E", X"3046", X"304E", 
X"3056", X"305F", X"3067", X"306F", X"3078", X"3080", X"3088", X"3090", X"3099", X"30A1", 
X"30A9", X"30B1", X"30BA", X"30C2", X"30CA", X"30D2", X"30DB", X"30E3", X"30EB", X"30F4", 
X"30FC", X"3104", X"310C", X"3115", X"311D", X"3125", X"312D", X"3136", X"313E", X"3146", 
X"314E", X"3157", X"315F", X"3167", X"316F", X"3178", X"3180", X"3188", X"3190", X"3198", 
X"31A1", X"31A9", X"31B1", X"31B9", X"31C2", X"31CA", X"31D2", X"31DA", X"31E3", X"31EB", 
X"31F3", X"31FB", X"3203", X"320C", X"3214", X"321C", X"3224", X"322D", X"3235", X"323D", 
X"3245", X"324D", X"3256", X"325E", X"3266", X"326E", X"3277", X"327F", X"3287", X"328F", 
X"3297", X"32A0", X"32A8", X"32B0", X"32B8", X"32C0", X"32C9", X"32D1", X"32D9", X"32E1", 
X"32E9", X"32F2", X"32FA", X"3302", X"330A", X"3312", X"331B", X"3323", X"332B", X"3333", 
X"333B", X"3344", X"334C", X"3354", X"335C", X"3364", X"336C", X"3375", X"337D", X"3385", 
X"338D", X"3395", X"339E", X"33A6", X"33AE", X"33B6", X"33BE", X"33C6", X"33CF", X"33D7", 
X"33DF", X"33E7", X"33EF", X"33F7", X"3400", X"3408", X"3410", X"3418", X"3420", X"3428", 
X"3431", X"3439", X"3441", X"3449", X"3451", X"3459", X"3462", X"346A", X"3472", X"347A", 
X"3482", X"348A", X"3492", X"349B", X"34A3", X"34AB", X"34B3", X"34BB", X"34C3", X"34CB", 
X"34D4", X"34DC", X"34E4", X"34EC", X"34F4", X"34FC", X"3504", X"350D", X"3515", X"351D", 
X"3525", X"352D", X"3535", X"353D", X"3545", X"354E", X"3556", X"355E", X"3566", X"356E", 
X"3576", X"357E", X"3586", X"358F", X"3597", X"359F", X"35A7", X"35AF", X"35B7", X"35BF", 
X"35C7", X"35CF", X"35D8", X"35E0", X"35E8", X"35F0", X"35F8", X"3600", X"3608", X"3610", 
X"3618", X"3620", X"3629", X"3631", X"3639", X"3641", X"3649", X"3651", X"3659", X"3661", 
X"3669", X"3671", X"3679", X"3682", X"368A", X"3692", X"369A", X"36A2", X"36AA", X"36B2", 
X"36BA", X"36C2", X"36CA", X"36D2", X"36DA", X"36E3", X"36EB", X"36F3", X"36FB", X"3703", 
X"370B", X"3713", X"371B", X"3723", X"372B", X"3733", X"373B", X"3743", X"374B", X"3753", 
X"375B", X"3764", X"376C", X"3774", X"377C", X"3784", X"378C", X"3794", X"379C", X"37A4", 
X"37AC", X"37B4", X"37BC", X"37C4", X"37CC", X"37D4", X"37DC", X"37E4", X"37EC", X"37F4", 
X"37FC", X"3804", X"380C", X"3815", X"381D", X"3825", X"382D", X"3835", X"383D", X"3845", 
X"384D", X"3855", X"385D", X"3865", X"386D", X"3875", X"387D", X"3885", X"388D", X"3895", 
X"389D", X"38A5", X"38AD", X"38B5", X"38BD", X"38C5", X"38CD", X"38D5", X"38DD", X"38E5", 
X"38ED", X"38F5", X"38FD", X"3905", X"390D", X"3915", X"391D", X"3925", X"392D", X"3935", 
X"393D", X"3945", X"394D", X"3955", X"395D", X"3965", X"396D", X"3975", X"397D", X"3985", 
X"398D", X"3995", X"399D", X"39A5", X"39AD", X"39B5", X"39BD", X"39C5", X"39CD", X"39D5", 
X"39DD", X"39E5", X"39ED", X"39F5", X"39FD", X"3A04", X"3A0C", X"3A14", X"3A1C", X"3A24", 
X"3A2C", X"3A34", X"3A3C", X"3A44", X"3A4C", X"3A54", X"3A5C", X"3A64", X"3A6C", X"3A74", 
X"3A7C", X"3A84", X"3A8C", X"3A94", X"3A9C", X"3AA4", X"3AAB", X"3AB3", X"3ABB", X"3AC3", 
X"3ACB", X"3AD3", X"3ADB", X"3AE3", X"3AEB", X"3AF3", X"3AFB", X"3B03", X"3B0B", X"3B13", 
X"3B1B", X"3B23", X"3B2A", X"3B32", X"3B3A", X"3B42", X"3B4A", X"3B52", X"3B5A", X"3B62", 
X"3B6A", X"3B72", X"3B7A", X"3B82", X"3B89", X"3B91", X"3B99", X"3BA1", X"3BA9", X"3BB1", 
X"3BB9", X"3BC1", X"3BC9", X"3BD1", X"3BD8", X"3BE0", X"3BE8", X"3BF0", X"3BF8", X"3C00", 
X"3C08", X"3C10", X"3C18", X"3C20", X"3C27", X"3C2F", X"3C37", X"3C3F", X"3C47", X"3C4F", 
X"3C57", X"3C5F", X"3C66", X"3C6E", X"3C76", X"3C7E", X"3C86", X"3C8E", X"3C96", X"3C9E", 
X"3CA5", X"3CAD", X"3CB5", X"3CBD", X"3CC5", X"3CCD", X"3CD5", X"3CDD", X"3CE4", X"3CEC", 
X"3CF4", X"3CFC", X"3D04", X"3D0C", X"3D14", X"3D1B", X"3D23", X"3D2B", X"3D33", X"3D3B", 
X"3D43", X"3D4A", X"3D52", X"3D5A", X"3D62", X"3D6A", X"3D72", X"3D7A", X"3D81", X"3D89", 
X"3D91", X"3D99", X"3DA1", X"3DA9", X"3DB0", X"3DB8", X"3DC0", X"3DC8", X"3DD0", X"3DD8", 
X"3DDF", X"3DE7", X"3DEF", X"3DF7", X"3DFF", X"3E06", X"3E0E", X"3E16", X"3E1E", X"3E26", 
X"3E2D", X"3E35", X"3E3D", X"3E45", X"3E4D", X"3E55", X"3E5C", X"3E64", X"3E6C", X"3E74", 
X"3E7C", X"3E83", X"3E8B", X"3E93", X"3E9B", X"3EA3", X"3EAA", X"3EB2", X"3EBA", X"3EC2", 
X"3EC9", X"3ED1", X"3ED9", X"3EE1", X"3EE9", X"3EF0", X"3EF8", X"3F00", X"3F08", X"3F10", 
X"3F17", X"3F1F", X"3F27", X"3F2F", X"3F36", X"3F3E", X"3F46", X"3F4E", X"3F55", X"3F5D", 
X"3F65", X"3F6D", X"3F75", X"3F7C", X"3F84", X"3F8C", X"3F94", X"3F9B", X"3FA3", X"3FAB", 
X"3FB3", X"3FBA", X"3FC2", X"3FCA", X"3FD2", X"3FD9", X"3FE1", X"3FE9", X"3FF1", X"3FF8", 
X"4000", X"4008", X"400F", X"4017", X"401F", X"4027", X"402E", X"4036", X"403E", X"4046", 
X"404D", X"4055", X"405D", X"4065", X"406C", X"4074", X"407C", X"4083", X"408B", X"4093", 
X"409B", X"40A2", X"40AA", X"40B2", X"40B9", X"40C1", X"40C9", X"40D1", X"40D8", X"40E0", 
X"40E8", X"40EF", X"40F7", X"40FF", X"4106", X"410E", X"4116", X"411E", X"4125", X"412D", 
X"4135", X"413C", X"4144", X"414C", X"4153", X"415B", X"4163", X"416A", X"4172", X"417A", 
X"4181", X"4189", X"4191", X"4198", X"41A0", X"41A8", X"41AF", X"41B7", X"41BF", X"41C6", 
X"41CE", X"41D6", X"41DD", X"41E5", X"41ED", X"41F4", X"41FC", X"4204", X"420B", X"4213", 
X"421B", X"4222", X"422A", X"4232", X"4239", X"4241", X"4249", X"4250", X"4258", X"4260", 
X"4267", X"426F", X"4276", X"427E", X"4286", X"428D", X"4295", X"429D", X"42A4", X"42AC", 
X"42B3", X"42BB", X"42C3", X"42CA", X"42D2", X"42DA", X"42E1", X"42E9", X"42F0", X"42F8", 
X"4300", X"4307", X"430F", X"4317", X"431E", X"4326", X"432D", X"4335", X"433D", X"4344", 
X"434C", X"4353", X"435B", X"4363", X"436A", X"4372", X"4379", X"4381", X"4389", X"4390", 
X"4398", X"439F", X"43A7", X"43AE", X"43B6", X"43BE", X"43C5", X"43CD", X"43D4", X"43DC", 
X"43E4", X"43EB", X"43F3", X"43FA", X"4402", X"4409", X"4411", X"4419", X"4420", X"4428", 
X"442F", X"4437", X"443E", X"4446", X"444D", X"4455", X"445D", X"4464", X"446C", X"4473", 
X"447B", X"4482", X"448A", X"4491", X"4499", X"44A1", X"44A8", X"44B0", X"44B7", X"44BF", 
X"44C6", X"44CE", X"44D5", X"44DD", X"44E4", X"44EC", X"44F3", X"44FB", X"4502", X"450A", 
X"4512", X"4519", X"4521", X"4528", X"4530", X"4537", X"453F", X"4546", X"454E", X"4555", 
X"455D", X"4564", X"456C", X"4573", X"457B", X"4582", X"458A", X"4591", X"4599", X"45A0", 
X"45A8", X"45AF", X"45B7", X"45BE", X"45C6", X"45CD", X"45D5", X"45DC", X"45E4", X"45EB", 
X"45F3", X"45FA", X"4602", X"4609", X"4611", X"4618", X"4620", X"4627", X"462E", X"4636", 
X"463D", X"4645", X"464C", X"4654", X"465B", X"4663", X"466A", X"4672", X"4679", X"4681", 
X"4688", X"4690", X"4697", X"469E", X"46A6", X"46AD", X"46B5", X"46BC", X"46C4", X"46CB", 
X"46D3", X"46DA", X"46E1", X"46E9", X"46F0", X"46F8", X"46FF", X"4707", X"470E", X"4715", 
X"471D", X"4724", X"472C", X"4733", X"473B", X"4742", X"4749", X"4751", X"4758", X"4760", 
X"4767", X"476F", X"4776", X"477D", X"4785", X"478C", X"4794", X"479B", X"47A2", X"47AA", 
X"47B1", X"47B9", X"47C0", X"47C7", X"47CF", X"47D6", X"47DE", X"47E5", X"47EC", X"47F4", 
X"47FB", X"4803", X"480A", X"4811", X"4819", X"4820", X"4828", X"482F", X"4836", X"483E", 
X"4845", X"484C", X"4854", X"485B", X"4863", X"486A", X"4871", X"4879", X"4880", X"4887", 
X"488F", X"4896", X"489D", X"48A5", X"48AC", X"48B4", X"48BB", X"48C2", X"48CA", X"48D1", 
X"48D8", X"48E0", X"48E7", X"48EE", X"48F6", X"48FD", X"4904", X"490C", X"4913", X"491A", 
X"4922", X"4929", X"4930", X"4938", X"493F", X"4946", X"494E", X"4955", X"495C", X"4964", 
X"496B", X"4972", X"497A", X"4981", X"4988", X"4990", X"4997", X"499E", X"49A5", X"49AD", 
X"49B4", X"49BB", X"49C3", X"49CA", X"49D1", X"49D9", X"49E0", X"49E7", X"49EE", X"49F6", 
X"49FD", X"4A04", X"4A0C", X"4A13", X"4A1A", X"4A22", X"4A29", X"4A30", X"4A37", X"4A3F", 
X"4A46", X"4A4D", X"4A54", X"4A5C", X"4A63", X"4A6A", X"4A72", X"4A79", X"4A80", X"4A87", 
X"4A8F", X"4A96", X"4A9D", X"4AA4", X"4AAC", X"4AB3", X"4ABA", X"4AC1", X"4AC9", X"4AD0", 
X"4AD7", X"4ADE", X"4AE6", X"4AED", X"4AF4", X"4AFB", X"4B03", X"4B0A", X"4B11", X"4B18", 
X"4B20", X"4B27", X"4B2E", X"4B35", X"4B3D", X"4B44", X"4B4B", X"4B52", X"4B59", X"4B61", 
X"4B68", X"4B6F", X"4B76", X"4B7E", X"4B85", X"4B8C", X"4B93", X"4B9A", X"4BA2", X"4BA9", 
X"4BB0", X"4BB7", X"4BBE", X"4BC6", X"4BCD", X"4BD4", X"4BDB", X"4BE2", X"4BEA", X"4BF1", 
X"4BF8", X"4BFF", X"4C06", X"4C0E", X"4C15", X"4C1C", X"4C23", X"4C2A", X"4C32", X"4C39", 
X"4C40", X"4C47", X"4C4E", X"4C55", X"4C5D", X"4C64", X"4C6B", X"4C72", X"4C79", X"4C80", 
X"4C88", X"4C8F", X"4C96", X"4C9D", X"4CA4", X"4CAB", X"4CB3", X"4CBA", X"4CC1", X"4CC8", 
X"4CCF", X"4CD6", X"4CDD", X"4CE5", X"4CEC", X"4CF3", X"4CFA", X"4D01", X"4D08", X"4D0F", 
X"4D17", X"4D1E", X"4D25", X"4D2C", X"4D33", X"4D3A", X"4D41", X"4D48", X"4D50", X"4D57", 
X"4D5E", X"4D65", X"4D6C", X"4D73", X"4D7A", X"4D81", X"4D88", X"4D90", X"4D97", X"4D9E", 
X"4DA5", X"4DAC", X"4DB3", X"4DBA", X"4DC1", X"4DC8", X"4DD0", X"4DD7", X"4DDE", X"4DE5", 
X"4DEC", X"4DF3", X"4DFA", X"4E01", X"4E08", X"4E0F", X"4E16", X"4E1D", X"4E25", X"4E2C", 
X"4E33", X"4E3A", X"4E41", X"4E48", X"4E4F", X"4E56", X"4E5D", X"4E64", X"4E6B", X"4E72", 
X"4E79", X"4E80", X"4E88", X"4E8F", X"4E96", X"4E9D", X"4EA4", X"4EAB", X"4EB2", X"4EB9", 
X"4EC0", X"4EC7", X"4ECE", X"4ED5", X"4EDC", X"4EE3", X"4EEA", X"4EF1", X"4EF8", X"4EFF", 
X"4F06", X"4F0D", X"4F14", X"4F1B", X"4F22", X"4F29", X"4F30", X"4F37", X"4F3E", X"4F45", 
X"4F4D", X"4F54", X"4F5B", X"4F62", X"4F69", X"4F70", X"4F77", X"4F7E", X"4F85", X"4F8C", 
X"4F93", X"4F9A", X"4FA1", X"4FA8", X"4FAF", X"4FB6", X"4FBD", X"4FC4", X"4FCB", X"4FD2", 
X"4FD8", X"4FDF", X"4FE6", X"4FED", X"4FF4", X"4FFB", X"5002", X"5009", X"5010", X"5017", 
X"501E", X"5025", X"502C", X"5033", X"503A", X"5041", X"5048", X"504F", X"5056", X"505D", 
X"5064", X"506B", X"5072", X"5079", X"5080", X"5087", X"508E", X"5095", X"509B", X"50A2", 
X"50A9", X"50B0", X"50B7", X"50BE", X"50C5", X"50CC", X"50D3", X"50DA", X"50E1", X"50E8", 
X"50EF", X"50F6", X"50FC", X"5103", X"510A", X"5111", X"5118", X"511F", X"5126", X"512D", 
X"5134", X"513B", X"5142", X"5149", X"514F", X"5156", X"515D", X"5164", X"516B", X"5172", 
X"5179", X"5180", X"5187", X"518D", X"5194", X"519B", X"51A2", X"51A9", X"51B0", X"51B7", 
X"51BE", X"51C5", X"51CB", X"51D2", X"51D9", X"51E0", X"51E7", X"51EE", X"51F5", X"51FB", 
X"5202", X"5209", X"5210", X"5217", X"521E", X"5225", X"522B", X"5232", X"5239", X"5240", 
X"5247", X"524E", X"5255", X"525B", X"5262", X"5269", X"5270", X"5277", X"527E", X"5284", 
X"528B", X"5292", X"5299", X"52A0", X"52A7", X"52AD", X"52B4", X"52BB", X"52C2", X"52C9", 
X"52CF", X"52D6", X"52DD", X"52E4", X"52EB", X"52F2", X"52F8", X"52FF", X"5306", X"530D", 
X"5314", X"531A", X"5321", X"5328", X"532F", X"5335", X"533C", X"5343", X"534A", X"5351", 
X"5357", X"535E", X"5365", X"536C", X"5373", X"5379", X"5380", X"5387", X"538E", X"5394", 
X"539B", X"53A2", X"53A9", X"53AF", X"53B6", X"53BD", X"53C4", X"53CA", X"53D1", X"53D8", 
X"53DF", X"53E6", X"53EC", X"53F3", X"53FA", X"5400", X"5407", X"540E", X"5415", X"541B", 
X"5422", X"5429", X"5430", X"5436", X"543D", X"5444", X"544B", X"5451", X"5458", X"545F", 
X"5465", X"546C", X"5473", X"547A", X"5480", X"5487", X"548E", X"5494", X"549B", X"54A2", 
X"54A9", X"54AF", X"54B6", X"54BD", X"54C3", X"54CA", X"54D1", X"54D7", X"54DE", X"54E5", 
X"54EB", X"54F2", X"54F9", X"5500", X"5506", X"550D", X"5514", X"551A", X"5521", X"5528", 
X"552E", X"5535", X"553C", X"5542", X"5549", X"5550", X"5556", X"555D", X"5564", X"556A", 
X"5571", X"5578", X"557E", X"5585", X"558B", X"5592", X"5599", X"559F", X"55A6", X"55AD", 
X"55B3", X"55BA", X"55C1", X"55C7", X"55CE", X"55D5", X"55DB", X"55E2", X"55E8", X"55EF", 
X"55F6", X"55FC", X"5603", X"560A", X"5610", X"5617", X"561D", X"5624", X"562B", X"5631", 
X"5638", X"563E", X"5645", X"564C", X"5652", X"5659", X"565F", X"5666", X"566D", X"5673", 
X"567A", X"5680", X"5687", X"568D", X"5694", X"569B", X"56A1", X"56A8", X"56AE", X"56B5", 
X"56BC", X"56C2", X"56C9", X"56CF", X"56D6", X"56DC", X"56E3", X"56EA", X"56F0", X"56F7", 
X"56FD", X"5704", X"570A", X"5711", X"5717", X"571E", X"5724", X"572B", X"5732", X"5738", 
X"573F", X"5745", X"574C", X"5752", X"5759", X"575F", X"5766", X"576C", X"5773", X"5779", 
X"5780", X"5786", X"578D", X"5794", X"579A", X"57A1", X"57A7", X"57AE", X"57B4", X"57BB", 
X"57C1", X"57C8", X"57CE", X"57D5", X"57DB", X"57E2", X"57E8", X"57EF", X"57F5", X"57FC", 
X"5802", X"5809", X"580F", X"5816", X"581C", X"5822", X"5829", X"582F", X"5836", X"583C", 
X"5843", X"5849", X"5850", X"5856", X"585D", X"5863", X"586A", X"5870", X"5877", X"587D", 
X"5884", X"588A", X"5890", X"5897", X"589D", X"58A4", X"58AA", X"58B1", X"58B7", X"58BE", 
X"58C4", X"58CA", X"58D1", X"58D7", X"58DE", X"58E4", X"58EB", X"58F1", X"58F7", X"58FE", 
X"5904", X"590B", X"5911", X"5918", X"591E", X"5924", X"592B", X"5931", X"5938", X"593E", 
X"5944", X"594B", X"5951", X"5958", X"595E", X"5964", X"596B", X"5971", X"5978", X"597E", 
X"5984", X"598B", X"5991", X"5998", X"599E", X"59A4", X"59AB", X"59B1", X"59B7", X"59BE", 
X"59C4", X"59CB", X"59D1", X"59D7", X"59DE", X"59E4", X"59EA", X"59F1", X"59F7", X"59FD", 
X"5A04", X"5A0A", X"5A10", X"5A17", X"5A1D", X"5A24", X"5A2A", X"5A30", X"5A37", X"5A3D", 
X"5A43", X"5A4A", X"5A50", X"5A56", X"5A5D", X"5A63", X"5A69", X"5A70", X"5A76", X"5A7C", 
X"5A82", X"5A89", X"5A8F", X"5A95", X"5A9C", X"5AA2", X"5AA8", X"5AAF", X"5AB5", X"5ABB", 
X"5AC2", X"5AC8", X"5ACE", X"5AD4", X"5ADB", X"5AE1", X"5AE7", X"5AEE", X"5AF4", X"5AFA", 
X"5B01", X"5B07", X"5B0D", X"5B13", X"5B1A", X"5B20", X"5B26", X"5B2C", X"5B33", X"5B39", 
X"5B3F", X"5B46", X"5B4C", X"5B52", X"5B58", X"5B5F", X"5B65", X"5B6B", X"5B71", X"5B78", 
X"5B7E", X"5B84", X"5B8A", X"5B91", X"5B97", X"5B9D", X"5BA3", X"5BAA", X"5BB0", X"5BB6", 
X"5BBC", X"5BC2", X"5BC9", X"5BCF", X"5BD5", X"5BDB", X"5BE2", X"5BE8", X"5BEE", X"5BF4", 
X"5BFA", X"5C01", X"5C07", X"5C0D", X"5C13", X"5C1A", X"5C20", X"5C26", X"5C2C", X"5C32", 
X"5C39", X"5C3F", X"5C45", X"5C4B", X"5C51", X"5C58", X"5C5E", X"5C64", X"5C6A", X"5C70", 
X"5C76", X"5C7D", X"5C83", X"5C89", X"5C8F", X"5C95", X"5C9B", X"5CA2", X"5CA8", X"5CAE", 
X"5CB4", X"5CBA", X"5CC0", X"5CC7", X"5CCD", X"5CD3", X"5CD9", X"5CDF", X"5CE5", X"5CEC", 
X"5CF2", X"5CF8", X"5CFE", X"5D04", X"5D0A", X"5D10", X"5D16", X"5D1D", X"5D23", X"5D29", 
X"5D2F", X"5D35", X"5D3B", X"5D41", X"5D48", X"5D4E", X"5D54", X"5D5A", X"5D60", X"5D66", 
X"5D6C", X"5D72", X"5D78", X"5D7F", X"5D85", X"5D8B", X"5D91", X"5D97", X"5D9D", X"5DA3", 
X"5DA9", X"5DAF", X"5DB5", X"5DBB", X"5DC2", X"5DC8", X"5DCE", X"5DD4", X"5DDA", X"5DE0", 
X"5DE6", X"5DEC", X"5DF2", X"5DF8", X"5DFE", X"5E04", X"5E0A", X"5E10", X"5E17", X"5E1D", 
X"5E23", X"5E29", X"5E2F", X"5E35", X"5E3B", X"5E41", X"5E47", X"5E4D", X"5E53", X"5E59", 
X"5E5F", X"5E65", X"5E6B", X"5E71", X"5E77", X"5E7D", X"5E83", X"5E89", X"5E8F", X"5E95", 
X"5E9B", X"5EA1", X"5EA7", X"5EAD", X"5EB3", X"5EB9", X"5EBF", X"5EC5", X"5ECB", X"5ED1", 
X"5ED7", X"5EDD", X"5EE3", X"5EE9", X"5EEF", X"5EF5", X"5EFB", X"5F01", X"5F07", X"5F0D", 
X"5F13", X"5F19", X"5F1F", X"5F25", X"5F2B", X"5F31", X"5F37", X"5F3D", X"5F43", X"5F49", 
X"5F4F", X"5F55", X"5F5B", X"5F61", X"5F67", X"5F6D", X"5F73", X"5F79", X"5F7F", X"5F85", 
X"5F8B", X"5F91", X"5F97", X"5F9D", X"5FA2", X"5FA8", X"5FAE", X"5FB4", X"5FBA", X"5FC0", 
X"5FC6", X"5FCC", X"5FD2", X"5FD8", X"5FDE", X"5FE4", X"5FEA", X"5FF0", X"5FF5", X"5FFB", 
X"6001", X"6007", X"600D", X"6013", X"6019", X"601F", X"6025", X"602B", X"6031", X"6036", 
X"603C", X"6042", X"6048", X"604E", X"6054", X"605A", X"6060", X"6065", X"606B", X"6071", 
X"6077", X"607D", X"6083", X"6089", X"608F", X"6094", X"609A", X"60A0", X"60A6", X"60AC", 
X"60B2", X"60B8", X"60BD", X"60C3", X"60C9", X"60CF", X"60D5", X"60DB", X"60E1", X"60E6", 
X"60EC", X"60F2", X"60F8", X"60FE", X"6104", X"6109", X"610F", X"6115", X"611B", X"6121", 
X"6126", X"612C", X"6132", X"6138", X"613E", X"6144", X"6149", X"614F", X"6155", X"615B", 
X"6161", X"6166", X"616C", X"6172", X"6178", X"617E", X"6183", X"6189", X"618F", X"6195", 
X"619A", X"61A0", X"61A6", X"61AC", X"61B2", X"61B7", X"61BD", X"61C3", X"61C9", X"61CE", 
X"61D4", X"61DA", X"61E0", X"61E5", X"61EB", X"61F1", X"61F7", X"61FD", X"6202", X"6208", 
X"620E", X"6213", X"6219", X"621F", X"6225", X"622A", X"6230", X"6236", X"623C", X"6241", 
X"6247", X"624D", X"6253", X"6258", X"625E", X"6264", X"6269", X"626F", X"6275", X"627B", 
X"6280", X"6286", X"628C", X"6291", X"6297", X"629D", X"62A2", X"62A8", X"62AE", X"62B4", 
X"62B9", X"62BF", X"62C5", X"62CA", X"62D0", X"62D6", X"62DB", X"62E1", X"62E7", X"62EC", 
X"62F2", X"62F8", X"62FD", X"6303", X"6309", X"630E", X"6314", X"631A", X"631F", X"6325", 
X"632B", X"6330", X"6336", X"633C", X"6341", X"6347", X"634C", X"6352", X"6358", X"635D", 
X"6363", X"6369", X"636E", X"6374", X"637A", X"637F", X"6385", X"638A", X"6390", X"6396", 
X"639B", X"63A1", X"63A6", X"63AC", X"63B2", X"63B7", X"63BD", X"63C2", X"63C8", X"63CE", 
X"63D3", X"63D9", X"63DE", X"63E4", X"63EA", X"63EF", X"63F5", X"63FA", X"6400", X"6406", 
X"640B", X"6411", X"6416", X"641C", X"6421", X"6427", X"642D", X"6432", X"6438", X"643D", 
X"6443", X"6448", X"644E", X"6453", X"6459", X"645E", X"6464", X"646A", X"646F", X"6475", 
X"647A", X"6480", X"6485", X"648B", X"6490", X"6496", X"649B", X"64A1", X"64A6", X"64AC", 
X"64B1", X"64B7", X"64BC", X"64C2", X"64C8", X"64CD", X"64D3", X"64D8", X"64DE", X"64E3", 
X"64E9", X"64EE", X"64F4", X"64F9", X"64FF", X"6504", X"6509", X"650F", X"6514", X"651A", 
X"651F", X"6525", X"652A", X"6530", X"6535", X"653B", X"6540", X"6546", X"654B", X"6551", 
X"6556", X"655C", X"6561", X"6566", X"656C", X"6571", X"6577", X"657C", X"6582", X"6587", 
X"658D", X"6592", X"6597", X"659D", X"65A2", X"65A8", X"65AD", X"65B3", X"65B8", X"65BD", 
X"65C3", X"65C8", X"65CE", X"65D3", X"65D9", X"65DE", X"65E3", X"65E9", X"65EE", X"65F4", 
X"65F9", X"65FE", X"6604", X"6609", X"660F", X"6614", X"6619", X"661F", X"6624", X"662A", 
X"662F", X"6634", X"663A", X"663F", X"6644", X"664A", X"664F", X"6655", X"665A", X"665F", 
X"6665", X"666A", X"666F", X"6675", X"667A", X"667F", X"6685", X"668A", X"668F", X"6695", 
X"669A", X"66A0", X"66A5", X"66AA", X"66B0", X"66B5", X"66BA", X"66C0", X"66C5", X"66CA", 
X"66D0", X"66D5", X"66DA", X"66DF", X"66E5", X"66EA", X"66EF", X"66F5", X"66FA", X"66FF", 
X"6705", X"670A", X"670F", X"6715", X"671A", X"671F", X"6724", X"672A", X"672F", X"6734", 
X"673A", X"673F", X"6744", X"6749", X"674F", X"6754", X"6759", X"675F", X"6764", X"6769", 
X"676E", X"6774", X"6779", X"677E", X"6783", X"6789", X"678E", X"6793", X"6798", X"679E", 
X"67A3", X"67A8", X"67AD", X"67B3", X"67B8", X"67BD", X"67C2", X"67C8", X"67CD", X"67D2", 
X"67D7", X"67DC", X"67E2", X"67E7", X"67EC", X"67F1", X"67F7", X"67FC", X"6801", X"6806", 
X"680B", X"6811", X"6816", X"681B", X"6820", X"6825", X"682B", X"6830", X"6835", X"683A", 
X"683F", X"6844", X"684A", X"684F", X"6854", X"6859", X"685E", X"6864", X"6869", X"686E", 
X"6873", X"6878", X"687D", X"6883", X"6888", X"688D", X"6892", X"6897", X"689C", X"68A1", 
X"68A7", X"68AC", X"68B1", X"68B6", X"68BB", X"68C0", X"68C5", X"68CB", X"68D0", X"68D5", 
X"68DA", X"68DF", X"68E4", X"68E9", X"68EE", X"68F4", X"68F9", X"68FE", X"6903", X"6908", 
X"690D", X"6912", X"6917", X"691C", X"6922", X"6927", X"692C", X"6931", X"6936", X"693B", 
X"6940", X"6945", X"694A", X"694F", X"6954", X"6959", X"695F", X"6964", X"6969", X"696E", 
X"6973", X"6978", X"697D", X"6982", X"6987", X"698C", X"6991", X"6996", X"699B", X"69A0", 
X"69A5", X"69AA", X"69AF", X"69B5", X"69BA", X"69BF", X"69C4", X"69C9", X"69CE", X"69D3", 
X"69D8", X"69DD", X"69E2", X"69E7", X"69EC", X"69F1", X"69F6", X"69FB", X"6A00", X"6A05", 
X"6A0A", X"6A0F", X"6A14", X"6A19", X"6A1E", X"6A23", X"6A28", X"6A2D", X"6A32", X"6A37", 
X"6A3C", X"6A41", X"6A46", X"6A4B", X"6A50", X"6A55", X"6A5A", X"6A5F", X"6A64", X"6A69", 
X"6A6E", X"6A73", X"6A78", X"6A7C", X"6A81", X"6A86", X"6A8B", X"6A90", X"6A95", X"6A9A", 
X"6A9F", X"6AA4", X"6AA9", X"6AAE", X"6AB3", X"6AB8", X"6ABD", X"6AC2", X"6AC7", X"6ACC", 
X"6AD0", X"6AD5", X"6ADA", X"6ADF", X"6AE4", X"6AE9", X"6AEE", X"6AF3", X"6AF8", X"6AFD", 
X"6B02", X"6B07", X"6B0B", X"6B10", X"6B15", X"6B1A", X"6B1F", X"6B24", X"6B29", X"6B2E", 
X"6B33", X"6B37", X"6B3C", X"6B41", X"6B46", X"6B4B", X"6B50", X"6B55", X"6B5A", X"6B5E", 
X"6B63", X"6B68", X"6B6D", X"6B72", X"6B77", X"6B7C", X"6B80", X"6B85", X"6B8A", X"6B8F", 
X"6B94", X"6B99", X"6B9D", X"6BA2", X"6BA7", X"6BAC", X"6BB1", X"6BB6", X"6BBA", X"6BBF", 
X"6BC4", X"6BC9", X"6BCE", X"6BD3", X"6BD7", X"6BDC", X"6BE1", X"6BE6", X"6BEB", X"6BEF", 
X"6BF4", X"6BF9", X"6BFE", X"6C03", X"6C07", X"6C0C", X"6C11", X"6C16", X"6C1B", X"6C1F", 
X"6C24", X"6C29", X"6C2E", X"6C32", X"6C37", X"6C3C", X"6C41", X"6C46", X"6C4A", X"6C4F", 
X"6C54", X"6C59", X"6C5D", X"6C62", X"6C67", X"6C6C", X"6C70", X"6C75", X"6C7A", X"6C7F", 
X"6C83", X"6C88", X"6C8D", X"6C92", X"6C96", X"6C9B", X"6CA0", X"6CA4", X"6CA9", X"6CAE", 
X"6CB3", X"6CB7", X"6CBC", X"6CC1", X"6CC6", X"6CCA", X"6CCF", X"6CD4", X"6CD8", X"6CDD", 
X"6CE2", X"6CE6", X"6CEB", X"6CF0", X"6CF5", X"6CF9", X"6CFE", X"6D03", X"6D07", X"6D0C", 
X"6D11", X"6D15", X"6D1A", X"6D1F", X"6D23", X"6D28", X"6D2D", X"6D31", X"6D36", X"6D3B", 
X"6D3F", X"6D44", X"6D49", X"6D4D", X"6D52", X"6D57", X"6D5B", X"6D60", X"6D64", X"6D69", 
X"6D6E", X"6D72", X"6D77", X"6D7C", X"6D80", X"6D85", X"6D8A", X"6D8E", X"6D93", X"6D97", 
X"6D9C", X"6DA1", X"6DA5", X"6DAA", X"6DAE", X"6DB3", X"6DB8", X"6DBC", X"6DC1", X"6DC5", 
X"6DCA", X"6DCF", X"6DD3", X"6DD8", X"6DDC", X"6DE1", X"6DE6", X"6DEA", X"6DEF", X"6DF3", 
X"6DF8", X"6DFC", X"6E01", X"6E06", X"6E0A", X"6E0F", X"6E13", X"6E18", X"6E1C", X"6E21", 
X"6E26", X"6E2A", X"6E2F", X"6E33", X"6E38", X"6E3C", X"6E41", X"6E45", X"6E4A", X"6E4E", 
X"6E53", X"6E57", X"6E5C", X"6E61", X"6E65", X"6E6A", X"6E6E", X"6E73", X"6E77", X"6E7C", 
X"6E80", X"6E85", X"6E89", X"6E8E", X"6E92", X"6E97", X"6E9B", X"6EA0", X"6EA4", X"6EA9", 
X"6EAD", X"6EB2", X"6EB6", X"6EBB", X"6EBF", X"6EC4", X"6EC8", X"6ECD", X"6ED1", X"6ED5", 
X"6EDA", X"6EDE", X"6EE3", X"6EE7", X"6EEC", X"6EF0", X"6EF5", X"6EF9", X"6EFE", X"6F02", 
X"6F06", X"6F0B", X"6F0F", X"6F14", X"6F18", X"6F1D", X"6F21", X"6F26", X"6F2A", X"6F2E", 
X"6F33", X"6F37", X"6F3C", X"6F40", X"6F45", X"6F49", X"6F4D", X"6F52", X"6F56", X"6F5B", 
X"6F5F", X"6F63", X"6F68", X"6F6C", X"6F71", X"6F75", X"6F79", X"6F7E", X"6F82", X"6F87", 
X"6F8B", X"6F8F", X"6F94", X"6F98", X"6F9C", X"6FA1", X"6FA5", X"6FAA", X"6FAE", X"6FB2", 
X"6FB7", X"6FBB", X"6FBF", X"6FC4", X"6FC8", X"6FCC", X"6FD1", X"6FD5", X"6FDA", X"6FDE", 
X"6FE2", X"6FE7", X"6FEB", X"6FEF", X"6FF4", X"6FF8", X"6FFC", X"7001", X"7005", X"7009", 
X"700D", X"7012", X"7016", X"701A", X"701F", X"7023", X"7027", X"702C", X"7030", X"7034", 
X"7039", X"703D", X"7041", X"7045", X"704A", X"704E", X"7052", X"7057", X"705B", X"705F", 
X"7063", X"7068", X"706C", X"7070", X"7075", X"7079", X"707D", X"7081", X"7086", X"708A", 
X"708E", X"7092", X"7097", X"709B", X"709F", X"70A3", X"70A8", X"70AC", X"70B0", X"70B4", 
X"70B9", X"70BD", X"70C1", X"70C5", X"70C9", X"70CE", X"70D2", X"70D6", X"70DA", X"70DF", 
X"70E3", X"70E7", X"70EB", X"70EF", X"70F4", X"70F8", X"70FC", X"7100", X"7104", X"7109", 
X"710D", X"7111", X"7115", X"7119", X"711E", X"7122", X"7126", X"712A", X"712E", X"7132", 
X"7137", X"713B", X"713F", X"7143", X"7147", X"714B", X"7150", X"7154", X"7158", X"715C", 
X"7160", X"7164", X"7168", X"716D", X"7171", X"7175", X"7179", X"717D", X"7181", X"7185", 
X"718A", X"718E", X"7192", X"7196", X"719A", X"719E", X"71A2", X"71A6", X"71AB", X"71AF", 
X"71B3", X"71B7", X"71BB", X"71BF", X"71C3", X"71C7", X"71CB", X"71CF", X"71D3", X"71D8", 
X"71DC", X"71E0", X"71E4", X"71E8", X"71EC", X"71F0", X"71F4", X"71F8", X"71FC", X"7200", 
X"7204", X"7208", X"720D", X"7211", X"7215", X"7219", X"721D", X"7221", X"7225", X"7229", 
X"722D", X"7231", X"7235", X"7239", X"723D", X"7241", X"7245", X"7249", X"724D", X"7251", 
X"7255", X"7259", X"725D", X"7261", X"7265", X"7269", X"726D", X"7271", X"7275", X"7279", 
X"727D", X"7281", X"7285", X"7289", X"728D", X"7291", X"7295", X"7299", X"729D", X"72A1", 
X"72A5", X"72A9", X"72AD", X"72B1", X"72B5", X"72B9", X"72BD", X"72C1", X"72C5", X"72C9", 
X"72CD", X"72D1", X"72D5", X"72D9", X"72DD", X"72E0", X"72E4", X"72E8", X"72EC", X"72F0", 
X"72F4", X"72F8", X"72FC", X"7300", X"7304", X"7308", X"730C", X"7310", X"7314", X"7317", 
X"731B", X"731F", X"7323", X"7327", X"732B", X"732F", X"7333", X"7337", X"733B", X"733E", 
X"7342", X"7346", X"734A", X"734E", X"7352", X"7356", X"735A", X"735D", X"7361", X"7365", 
X"7369", X"736D", X"7371", X"7375", X"7379", X"737C", X"7380", X"7384", X"7388", X"738C", 
X"7390", X"7393", X"7397", X"739B", X"739F", X"73A3", X"73A7", X"73AA", X"73AE", X"73B2", 
X"73B6", X"73BA", X"73BE", X"73C1", X"73C5", X"73C9", X"73CD", X"73D1", X"73D4", X"73D8", 
X"73DC", X"73E0", X"73E4", X"73E7", X"73EB", X"73EF", X"73F3", X"73F7", X"73FA", X"73FE", 
X"7402", X"7406", X"7409", X"740D", X"7411", X"7415", X"7419", X"741C", X"7420", X"7424", 
X"7428", X"742B", X"742F", X"7433", X"7437", X"743A", X"743E", X"7442", X"7446", X"7449", 
X"744D", X"7451", X"7454", X"7458", X"745C", X"7460", X"7463", X"7467", X"746B", X"746E", 
X"7472", X"7476", X"747A", X"747D", X"7481", X"7485", X"7488", X"748C", X"7490", X"7493", 
X"7497", X"749B", X"749F", X"74A2", X"74A6", X"74AA", X"74AD", X"74B1", X"74B5", X"74B8", 
X"74BC", X"74C0", X"74C3", X"74C7", X"74CB", X"74CE", X"74D2", X"74D6", X"74D9", X"74DD", 
X"74E1", X"74E4", X"74E8", X"74EB", X"74EF", X"74F3", X"74F6", X"74FA", X"74FE", X"7501", 
X"7505", X"7508", X"750C", X"7510", X"7513", X"7517", X"751B", X"751E", X"7522", X"7525", 
X"7529", X"752D", X"7530", X"7534", X"7537", X"753B", X"753E", X"7542", X"7546", X"7549", 
X"754D", X"7550", X"7554", X"7558", X"755B", X"755F", X"7562", X"7566", X"7569", X"756D", 
X"7570", X"7574", X"7578", X"757B", X"757F", X"7582", X"7586", X"7589", X"758D", X"7590", 
X"7594", X"7597", X"759B", X"759E", X"75A2", X"75A6", X"75A9", X"75AD", X"75B0", X"75B4", 
X"75B7", X"75BB", X"75BE", X"75C2", X"75C5", X"75C9", X"75CC", X"75D0", X"75D3", X"75D7", 
X"75DA", X"75DE", X"75E1", X"75E5", X"75E8", X"75EB", X"75EF", X"75F2", X"75F6", X"75F9", 
X"75FD", X"7600", X"7604", X"7607", X"760B", X"760E", X"7612", X"7615", X"7618", X"761C", 
X"761F", X"7623", X"7626", X"762A", X"762D", X"7631", X"7634", X"7637", X"763B", X"763E", 
X"7642", X"7645", X"7649", X"764C", X"764F", X"7653", X"7656", X"765A", X"765D", X"7660", 
X"7664", X"7667", X"766B", X"766E", X"7671", X"7675", X"7678", X"767B", X"767F", X"7682", 
X"7686", X"7689", X"768C", X"7690", X"7693", X"7696", X"769A", X"769D", X"76A1", X"76A4", 
X"76A7", X"76AB", X"76AE", X"76B1", X"76B5", X"76B8", X"76BB", X"76BF", X"76C2", X"76C5", 
X"76C9", X"76CC", X"76CF", X"76D3", X"76D6", X"76D9", X"76DD", X"76E0", X"76E3", X"76E7", 
X"76EA", X"76ED", X"76F0", X"76F4", X"76F7", X"76FA", X"76FE", X"7701", X"7704", X"7708", 
X"770B", X"770E", X"7711", X"7715", X"7718", X"771B", X"771E", X"7722", X"7725", X"7728", 
X"772C", X"772F", X"7732", X"7735", X"7739", X"773C", X"773F", X"7742", X"7746", X"7749", 
X"774C", X"774F", X"7753", X"7756", X"7759", X"775C", X"775F", X"7763", X"7766", X"7769", 
X"776C", X"7770", X"7773", X"7776", X"7779", X"777C", X"7780", X"7783", X"7786", X"7789", 
X"778C", X"7790", X"7793", X"7796", X"7799", X"779C", X"779F", X"77A3", X"77A6", X"77A9", 
X"77AC", X"77AF", X"77B3", X"77B6", X"77B9", X"77BC", X"77BF", X"77C2", X"77C5", X"77C9", 
X"77CC", X"77CF", X"77D2", X"77D5", X"77D8", X"77DB", X"77DF", X"77E2", X"77E5", X"77E8", 
X"77EB", X"77EE", X"77F1", X"77F4", X"77F8", X"77FB", X"77FE", X"7801", X"7804", X"7807", 
X"780A", X"780D", X"7810", X"7814", X"7817", X"781A", X"781D", X"7820", X"7823", X"7826", 
X"7829", X"782C", X"782F", X"7832", X"7835", X"7839", X"783C", X"783F", X"7842", X"7845", 
X"7848", X"784B", X"784E", X"7851", X"7854", X"7857", X"785A", X"785D", X"7860", X"7863", 
X"7866", X"7869", X"786C", X"786F", X"7872", X"7875", X"7878", X"787B", X"787E", X"7882", 
X"7885", X"7888", X"788B", X"788E", X"7891", X"7894", X"7897", X"789A", X"789D", X"78A0", 
X"78A3", X"78A5", X"78A8", X"78AB", X"78AE", X"78B1", X"78B4", X"78B7", X"78BA", X"78BD", 
X"78C0", X"78C3", X"78C6", X"78C9", X"78CC", X"78CF", X"78D2", X"78D5", X"78D8", X"78DB", 
X"78DE", X"78E1", X"78E4", X"78E7", X"78EA", X"78EC", X"78EF", X"78F2", X"78F5", X"78F8", 
X"78FB", X"78FE", X"7901", X"7904", X"7907", X"790A", X"790D", X"790F", X"7912", X"7915", 
X"7918", X"791B", X"791E", X"7921", X"7924", X"7927", X"7929", X"792C", X"792F", X"7932", 
X"7935", X"7938", X"793B", X"793E", X"7940", X"7943", X"7946", X"7949", X"794C", X"794F", 
X"7952", X"7954", X"7957", X"795A", X"795D", X"7960", X"7963", X"7966", X"7968", X"796B", 
X"796E", X"7971", X"7974", X"7976", X"7979", X"797C", X"797F", X"7982", X"7985", X"7987", 
X"798A", X"798D", X"7990", X"7993", X"7995", X"7998", X"799B", X"799E", X"79A0", X"79A3", 
X"79A6", X"79A9", X"79AC", X"79AE", X"79B1", X"79B4", X"79B7", X"79B9", X"79BC", X"79BF", 
X"79C2", X"79C4", X"79C7", X"79CA", X"79CD", X"79CF", X"79D2", X"79D5", X"79D8", X"79DA", 
X"79DD", X"79E0", X"79E3", X"79E5", X"79E8", X"79EB", X"79EE", X"79F0", X"79F3", X"79F6", 
X"79F8", X"79FB", X"79FE", X"7A01", X"7A03", X"7A06", X"7A09", X"7A0B", X"7A0E", X"7A11", 
X"7A13", X"7A16", X"7A19", X"7A1B", X"7A1E", X"7A21", X"7A23", X"7A26", X"7A29", X"7A2B", 
X"7A2E", X"7A31", X"7A33", X"7A36", X"7A39", X"7A3B", X"7A3E", X"7A41", X"7A43", X"7A46", 
X"7A49", X"7A4B", X"7A4E", X"7A51", X"7A53", X"7A56", X"7A58", X"7A5B", X"7A5E", X"7A60", 
X"7A63", X"7A66", X"7A68", X"7A6B", X"7A6D", X"7A70", X"7A73", X"7A75", X"7A78", X"7A7A", 
X"7A7D", X"7A80", X"7A82", X"7A85", X"7A87", X"7A8A", X"7A8D", X"7A8F", X"7A92", X"7A94", 
X"7A97", X"7A99", X"7A9C", X"7A9F", X"7AA1", X"7AA4", X"7AA6", X"7AA9", X"7AAB", X"7AAE", 
X"7AB0", X"7AB3", X"7AB6", X"7AB8", X"7ABB", X"7ABD", X"7AC0", X"7AC2", X"7AC5", X"7AC7", 
X"7ACA", X"7ACC", X"7ACF", X"7AD1", X"7AD4", X"7AD6", X"7AD9", X"7ADB", X"7ADE", X"7AE0", 
X"7AE3", X"7AE5", X"7AE8", X"7AEA", X"7AED", X"7AEF", X"7AF2", X"7AF4", X"7AF7", X"7AF9", 
X"7AFC", X"7AFE", X"7B01", X"7B03", X"7B06", X"7B08", X"7B0B", X"7B0D", X"7B10", X"7B12", 
X"7B14", X"7B17", X"7B19", X"7B1C", X"7B1E", X"7B21", X"7B23", X"7B26", X"7B28", X"7B2A", 
X"7B2D", X"7B2F", X"7B32", X"7B34", X"7B37", X"7B39", X"7B3B", X"7B3E", X"7B40", X"7B43", 
X"7B45", X"7B47", X"7B4A", X"7B4C", X"7B4F", X"7B51", X"7B53", X"7B56", X"7B58", X"7B5B", 
X"7B5D", X"7B5F", X"7B62", X"7B64", X"7B67", X"7B69", X"7B6B", X"7B6E", X"7B70", X"7B72", 
X"7B75", X"7B77", X"7B79", X"7B7C", X"7B7E", X"7B81", X"7B83", X"7B85", X"7B88", X"7B8A", 
X"7B8C", X"7B8F", X"7B91", X"7B93", X"7B96", X"7B98", X"7B9A", X"7B9D", X"7B9F", X"7BA1", 
X"7BA3", X"7BA6", X"7BA8", X"7BAA", X"7BAD", X"7BAF", X"7BB1", X"7BB4", X"7BB6", X"7BB8", 
X"7BBA", X"7BBD", X"7BBF", X"7BC1", X"7BC4", X"7BC6", X"7BC8", X"7BCA", X"7BCD", X"7BCF", 
X"7BD1", X"7BD4", X"7BD6", X"7BD8", X"7BDA", X"7BDD", X"7BDF", X"7BE1", X"7BE3", X"7BE6", 
X"7BE8", X"7BEA", X"7BEC", X"7BEE", X"7BF1", X"7BF3", X"7BF5", X"7BF7", X"7BFA", X"7BFC", 
X"7BFE", X"7C00", X"7C03", X"7C05", X"7C07", X"7C09", X"7C0B", X"7C0E", X"7C10", X"7C12", 
X"7C14", X"7C16", X"7C19", X"7C1B", X"7C1D", X"7C1F", X"7C21", X"7C23", X"7C26", X"7C28", 
X"7C2A", X"7C2C", X"7C2E", X"7C30", X"7C33", X"7C35", X"7C37", X"7C39", X"7C3B", X"7C3D", 
X"7C40", X"7C42", X"7C44", X"7C46", X"7C48", X"7C4A", X"7C4C", X"7C4F", X"7C51", X"7C53", 
X"7C55", X"7C57", X"7C59", X"7C5B", X"7C5D", X"7C60", X"7C62", X"7C64", X"7C66", X"7C68", 
X"7C6A", X"7C6C", X"7C6E", X"7C70", X"7C72", X"7C75", X"7C77", X"7C79", X"7C7B", X"7C7D", 
X"7C7F", X"7C81", X"7C83", X"7C85", X"7C87", X"7C89", X"7C8B", X"7C8D", X"7C8F", X"7C92", 
X"7C94", X"7C96", X"7C98", X"7C9A", X"7C9C", X"7C9E", X"7CA0", X"7CA2", X"7CA4", X"7CA6", 
X"7CA8", X"7CAA", X"7CAC", X"7CAE", X"7CB0", X"7CB2", X"7CB4", X"7CB6", X"7CB8", X"7CBA", 
X"7CBC", X"7CBE", X"7CC0", X"7CC2", X"7CC4", X"7CC6", X"7CC8", X"7CCA", X"7CCC", X"7CCE", 
X"7CD0", X"7CD2", X"7CD4", X"7CD6", X"7CD8", X"7CDA", X"7CDC", X"7CDE", X"7CE0", X"7CE2", 
X"7CE4", X"7CE6", X"7CE8", X"7CEA", X"7CEC", X"7CEE", X"7CF0", X"7CF1", X"7CF3", X"7CF5", 
X"7CF7", X"7CF9", X"7CFB", X"7CFD", X"7CFF", X"7D01", X"7D03", X"7D05", X"7D07", X"7D09", 
X"7D0A", X"7D0C", X"7D0E", X"7D10", X"7D12", X"7D14", X"7D16", X"7D18", X"7D1A", X"7D1C", 
X"7D1D", X"7D1F", X"7D21", X"7D23", X"7D25", X"7D27", X"7D29", X"7D2B", X"7D2C", X"7D2E", 
X"7D30", X"7D32", X"7D34", X"7D36", X"7D38", X"7D3A", X"7D3B", X"7D3D", X"7D3F", X"7D41", 
X"7D43", X"7D45", X"7D46", X"7D48", X"7D4A", X"7D4C", X"7D4E", X"7D50", X"7D51", X"7D53", 
X"7D55", X"7D57", X"7D59", X"7D5A", X"7D5C", X"7D5E", X"7D60", X"7D62", X"7D63", X"7D65", 
X"7D67", X"7D69", X"7D6B", X"7D6C", X"7D6E", X"7D70", X"7D72", X"7D74", X"7D75", X"7D77", 
X"7D79", X"7D7B", X"7D7C", X"7D7E", X"7D80", X"7D82", X"7D83", X"7D85", X"7D87", X"7D89", 
X"7D8A", X"7D8C", X"7D8E", X"7D90", X"7D91", X"7D93", X"7D95", X"7D97", X"7D98", X"7D9A", 
X"7D9C", X"7D9D", X"7D9F", X"7DA1", X"7DA3", X"7DA4", X"7DA6", X"7DA8", X"7DA9", X"7DAB", 
X"7DAD", X"7DAE", X"7DB0", X"7DB2", X"7DB4", X"7DB5", X"7DB7", X"7DB9", X"7DBA", X"7DBC", 
X"7DBE", X"7DBF", X"7DC1", X"7DC3", X"7DC4", X"7DC6", X"7DC8", X"7DC9", X"7DCB", X"7DCD", 
X"7DCE", X"7DD0", X"7DD1", X"7DD3", X"7DD5", X"7DD6", X"7DD8", X"7DDA", X"7DDB", X"7DDD", 
X"7DDF", X"7DE0", X"7DE2", X"7DE3", X"7DE5", X"7DE7", X"7DE8", X"7DEA", X"7DEB", X"7DED", 
X"7DEF", X"7DF0", X"7DF2", X"7DF3", X"7DF5", X"7DF7", X"7DF8", X"7DFA", X"7DFB", X"7DFD", 
X"7DFF", X"7E00", X"7E02", X"7E03", X"7E05", X"7E06", X"7E08", X"7E0A", X"7E0B", X"7E0D", 
X"7E0E", X"7E10", X"7E11", X"7E13", X"7E14", X"7E16", X"7E17", X"7E19", X"7E1B", X"7E1C", 
X"7E1E", X"7E1F", X"7E21", X"7E22", X"7E24", X"7E25", X"7E27", X"7E28", X"7E2A", X"7E2B", 
X"7E2D", X"7E2E", X"7E30", X"7E31", X"7E33", X"7E34", X"7E36", X"7E37", X"7E39", X"7E3A", 
X"7E3C", X"7E3D", X"7E3F", X"7E40", X"7E42", X"7E43", X"7E44", X"7E46", X"7E47", X"7E49", 
X"7E4A", X"7E4C", X"7E4D", X"7E4F", X"7E50", X"7E52", X"7E53", X"7E54", X"7E56", X"7E57", 
X"7E59", X"7E5A", X"7E5C", X"7E5D", X"7E5E", X"7E60", X"7E61", X"7E63", X"7E64", X"7E66", 
X"7E67", X"7E68", X"7E6A", X"7E6B", X"7E6D", X"7E6E", X"7E6F", X"7E71", X"7E72", X"7E74", 
X"7E75", X"7E76", X"7E78", X"7E79", X"7E7A", X"7E7C", X"7E7D", X"7E7F", X"7E80", X"7E81", 
X"7E83", X"7E84", X"7E85", X"7E87", X"7E88", X"7E89", X"7E8B", X"7E8C", X"7E8D", X"7E8F", 
X"7E90", X"7E91", X"7E93", X"7E94", X"7E95", X"7E97", X"7E98", X"7E99", X"7E9B", X"7E9C", 
X"7E9D", X"7E9F", X"7EA0", X"7EA1", X"7EA3", X"7EA4", X"7EA5", X"7EA6", X"7EA8", X"7EA9", 
X"7EAA", X"7EAC", X"7EAD", X"7EAE", X"7EAF", X"7EB1", X"7EB2", X"7EB3", X"7EB5", X"7EB6", 
X"7EB7", X"7EB8", X"7EBA", X"7EBB", X"7EBC", X"7EBD", X"7EBF", X"7EC0", X"7EC1", X"7EC2", 
X"7EC4", X"7EC5", X"7EC6", X"7EC7", X"7EC9", X"7ECA", X"7ECB", X"7ECC", X"7ECD", X"7ECF", 
X"7ED0", X"7ED1", X"7ED2", X"7ED3", X"7ED5", X"7ED6", X"7ED7", X"7ED8", X"7ED9", X"7EDB", 
X"7EDC", X"7EDD", X"7EDE", X"7EDF", X"7EE1", X"7EE2", X"7EE3", X"7EE4", X"7EE5", X"7EE6", 
X"7EE8", X"7EE9", X"7EEA", X"7EEB", X"7EEC", X"7EED", X"7EEF", X"7EF0", X"7EF1", X"7EF2", 
X"7EF3", X"7EF4", X"7EF5", X"7EF7", X"7EF8", X"7EF9", X"7EFA", X"7EFB", X"7EFC", X"7EFD", 
X"7EFF", X"7F00", X"7F01", X"7F02", X"7F03", X"7F04", X"7F05", X"7F06", X"7F07", X"7F08", 
X"7F0A", X"7F0B", X"7F0C", X"7F0D", X"7F0E", X"7F0F", X"7F10", X"7F11", X"7F12", X"7F13", 
X"7F14", X"7F15", X"7F17", X"7F18", X"7F19", X"7F1A", X"7F1B", X"7F1C", X"7F1D", X"7F1E", 
X"7F1F", X"7F20", X"7F21", X"7F22", X"7F23", X"7F24", X"7F25", X"7F26", X"7F27", X"7F28", 
X"7F29", X"7F2A", X"7F2B", X"7F2C", X"7F2D", X"7F2E", X"7F2F", X"7F30", X"7F31", X"7F32", 
X"7F33", X"7F34", X"7F35", X"7F36", X"7F37", X"7F38", X"7F39", X"7F3A", X"7F3B", X"7F3C", 
X"7F3D", X"7F3E", X"7F3F", X"7F40", X"7F41", X"7F42", X"7F43", X"7F44", X"7F45", X"7F46", 
X"7F47", X"7F48", X"7F49", X"7F4A", X"7F4B", X"7F4C", X"7F4C", X"7F4D", X"7F4E", X"7F4F", 
X"7F50", X"7F51", X"7F52", X"7F53", X"7F54", X"7F55", X"7F56", X"7F57", X"7F58", X"7F58", 
X"7F59", X"7F5A", X"7F5B", X"7F5C", X"7F5D", X"7F5E", X"7F5F", X"7F60", X"7F60", X"7F61", 
X"7F62", X"7F63", X"7F64", X"7F65", X"7F66", X"7F67", X"7F67", X"7F68", X"7F69", X"7F6A", 
X"7F6B", X"7F6C", X"7F6D", X"7F6D", X"7F6E", X"7F6F", X"7F70", X"7F71", X"7F72", X"7F72", 
X"7F73", X"7F74", X"7F75", X"7F76", X"7F77", X"7F77", X"7F78", X"7F79", X"7F7A", X"7F7B", 
X"7F7B", X"7F7C", X"7F7D", X"7F7E", X"7F7F", X"7F7F", X"7F80", X"7F81", X"7F82", X"7F83", 
X"7F83", X"7F84", X"7F85", X"7F86", X"7F86", X"7F87", X"7F88", X"7F89", X"7F89", X"7F8A", 
X"7F8B", X"7F8C", X"7F8C", X"7F8D", X"7F8E", X"7F8F", X"7F8F", X"7F90", X"7F91", X"7F92", 
X"7F92", X"7F93", X"7F94", X"7F95", X"7F95", X"7F96", X"7F97", X"7F97", X"7F98", X"7F99", 
X"7F9A", X"7F9A", X"7F9B", X"7F9C", X"7F9C", X"7F9D", X"7F9E", X"7F9E", X"7F9F", X"7FA0", 
X"7FA1", X"7FA1", X"7FA2", X"7FA3", X"7FA3", X"7FA4", X"7FA5", X"7FA5", X"7FA6", X"7FA7", 
X"7FA7", X"7FA8", X"7FA9", X"7FA9", X"7FAA", X"7FAA", X"7FAB", X"7FAC", X"7FAC", X"7FAD", 
X"7FAE", X"7FAE", X"7FAF", X"7FB0", X"7FB0", X"7FB1", X"7FB1", X"7FB2", X"7FB3", X"7FB3", 
X"7FB4", X"7FB4", X"7FB5", X"7FB6", X"7FB6", X"7FB7", X"7FB7", X"7FB8", X"7FB9", X"7FB9", 
X"7FBA", X"7FBA", X"7FBB", X"7FBC", X"7FBC", X"7FBD", X"7FBD", X"7FBE", X"7FBE", X"7FBF", 
X"7FC0", X"7FC0", X"7FC1", X"7FC1", X"7FC2", X"7FC2", X"7FC3", X"7FC3", X"7FC4", X"7FC5", 
X"7FC5", X"7FC6", X"7FC6", X"7FC7", X"7FC7", X"7FC8", X"7FC8", X"7FC9", X"7FC9", X"7FCA", 
X"7FCA", X"7FCB", X"7FCB", X"7FCC", X"7FCC", X"7FCD", X"7FCD", X"7FCE", X"7FCE", X"7FCF", 
X"7FCF", X"7FD0", X"7FD0", X"7FD1", X"7FD1", X"7FD2", X"7FD2", X"7FD3", X"7FD3", X"7FD4", 
X"7FD4", X"7FD4", X"7FD5", X"7FD5", X"7FD6", X"7FD6", X"7FD7", X"7FD7", X"7FD8", X"7FD8", 
X"7FD9", X"7FD9", X"7FD9", X"7FDA", X"7FDA", X"7FDB", X"7FDB", X"7FDC", X"7FDC", X"7FDC", 
X"7FDD", X"7FDD", X"7FDE", X"7FDE", X"7FDE", X"7FDF", X"7FDF", X"7FE0", X"7FE0", X"7FE0", 
X"7FE1", X"7FE1", X"7FE2", X"7FE2", X"7FE2", X"7FE3", X"7FE3", X"7FE3", X"7FE4", X"7FE4", 
X"7FE5", X"7FE5", X"7FE5", X"7FE6", X"7FE6", X"7FE6", X"7FE7", X"7FE7", X"7FE7", X"7FE8", 
X"7FE8", X"7FE8", X"7FE9", X"7FE9", X"7FE9", X"7FEA", X"7FEA", X"7FEA", X"7FEB", X"7FEB", 
X"7FEB", X"7FEC", X"7FEC", X"7FEC", X"7FED", X"7FED", X"7FED", X"7FEE", X"7FEE", X"7FEE", 
X"7FEE", X"7FEF", X"7FEF", X"7FEF", X"7FF0", X"7FF0", X"7FF0", X"7FF0", X"7FF1", X"7FF1", 
X"7FF1", X"7FF2", X"7FF2", X"7FF2", X"7FF2", X"7FF3", X"7FF3", X"7FF3", X"7FF3", X"7FF4", 
X"7FF4", X"7FF4", X"7FF4", X"7FF5", X"7FF5", X"7FF5", X"7FF5", X"7FF5", X"7FF6", X"7FF6", 
X"7FF6", X"7FF6", X"7FF7", X"7FF7", X"7FF7", X"7FF7", X"7FF7", X"7FF8", X"7FF8", X"7FF8", 
X"7FF8", X"7FF8", X"7FF9", X"7FF9", X"7FF9", X"7FF9", X"7FF9", X"7FFA", X"7FFA", X"7FFA", 
X"7FFA", X"7FFA", X"7FFA", X"7FFB", X"7FFB", X"7FFB", X"7FFB", X"7FFB", X"7FFB", X"7FFB", 
X"7FFC", X"7FFC", X"7FFC", X"7FFC", X"7FFC", X"7FFC", X"7FFC", X"7FFD", X"7FFD", X"7FFD", 
X"7FFD", X"7FFD", X"7FFD", X"7FFD", X"7FFD", X"7FFE", X"7FFE", X"7FFE", X"7FFE", X"7FFE", 
X"7FFE", X"7FFE", X"7FFE", X"7FFE", X"7FFE", X"7FFF", X"7FFF", X"7FFF", X"7FFF", X"7FFF", 
X"7FFF", X"7FFF", X"7FFF", X"7FFF", X"7FFF", X"7FFF", X"7FFF", X"7FFF", X"7FFF", X"7FFF", 
X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", 
X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000", X"8000"
);
begin
	process(H)
	begin
		if(H'event and H='1')then
			COSINUS <= TABLE(TO_INTEGER(UNSIGNED(ANGLE)));
		end if;
	end process;
end architecture;